VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_carry_ripple_7_bit
  CLASS BLOCK ;
  FOREIGN tt_um_carry_ripple_7_bit ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.621000 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.335899 ;
    ANTENNADIFFAREA 18.907700 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.800500 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.800500 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.800500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.800500 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.800500 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.800500 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.800500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 30.600 202.650 78.700 204.310 ;
      LAYER pwell ;
        RECT 32.950 202.365 33.350 202.400 ;
        RECT 36.300 202.365 37.150 202.450 ;
        RECT 39.000 202.365 39.500 202.400 ;
        RECT 42.500 202.365 44.350 202.400 ;
        RECT 45.500 202.365 47.100 202.450 ;
        RECT 50.050 202.365 50.900 202.400 ;
        RECT 52.750 202.365 53.600 202.400 ;
        RECT 56.550 202.365 58.450 202.400 ;
        RECT 60.050 202.365 61.150 202.400 ;
        RECT 64.100 202.365 65.000 202.400 ;
        RECT 66.600 202.365 67.700 202.450 ;
        RECT 70.650 202.365 72.600 202.400 ;
        RECT 74.250 202.365 75.400 202.450 ;
        RECT 31.945 202.275 32.895 202.365 ;
        RECT 30.965 201.455 32.895 202.275 ;
        RECT 32.950 202.275 37.150 202.365 ;
        RECT 38.015 202.275 38.965 202.365 ;
        RECT 32.950 201.550 38.965 202.275 ;
        RECT 33.245 201.500 38.965 201.550 ;
        RECT 39.000 202.275 44.350 202.365 ;
        RECT 45.235 202.275 50.900 202.365 ;
        RECT 51.785 202.275 52.735 202.365 ;
        RECT 39.000 201.500 52.735 202.275 ;
        RECT 52.750 202.275 58.450 202.365 ;
        RECT 59.335 202.275 65.000 202.365 ;
        RECT 65.885 202.275 72.600 202.365 ;
        RECT 73.495 202.275 78.465 202.365 ;
        RECT 52.750 201.500 78.465 202.275 ;
        RECT 33.245 201.455 36.975 201.500 ;
        RECT 30.965 201.435 31.115 201.455 ;
        RECT 30.945 201.265 31.115 201.435 ;
        RECT 33.345 201.265 33.515 201.455 ;
        RECT 36.345 201.105 36.975 201.455 ;
        RECT 37.035 201.455 38.965 201.500 ;
        RECT 37.035 201.435 37.185 201.455 ;
        RECT 37.015 201.265 37.185 201.435 ;
        RECT 39.125 201.110 39.400 201.500 ;
        RECT 39.415 201.455 42.585 201.500 ;
        RECT 44.255 201.455 46.185 201.500 ;
        RECT 46.985 201.455 50.155 201.500 ;
        RECT 50.805 201.455 52.735 201.500 ;
        RECT 53.485 201.455 56.655 201.500 ;
        RECT 58.355 201.455 60.285 201.500 ;
        RECT 61.035 201.455 64.205 201.500 ;
        RECT 64.905 201.455 66.835 201.500 ;
        RECT 67.585 201.455 70.755 201.500 ;
        RECT 72.515 201.455 74.445 201.500 ;
        RECT 75.295 201.455 78.465 201.500 ;
        RECT 39.515 201.265 39.685 201.455 ;
        RECT 44.255 201.435 44.405 201.455 ;
        RECT 44.235 201.265 44.405 201.435 ;
        RECT 47.085 201.265 47.255 201.455 ;
        RECT 50.805 201.435 50.955 201.455 ;
        RECT 50.785 201.265 50.955 201.435 ;
        RECT 53.585 201.265 53.755 201.455 ;
        RECT 58.355 201.435 58.505 201.455 ;
        RECT 58.335 201.265 58.505 201.435 ;
        RECT 61.135 201.265 61.305 201.455 ;
        RECT 64.905 201.435 65.055 201.455 ;
        RECT 64.885 201.265 65.055 201.435 ;
        RECT 67.685 201.265 67.855 201.455 ;
        RECT 72.515 201.435 72.665 201.455 ;
        RECT 72.495 201.265 72.665 201.435 ;
        RECT 75.395 201.265 75.565 201.455 ;
      LAYER nwell ;
        RECT 43.500 200.910 44.350 200.960 ;
        RECT 71.800 200.920 72.650 200.950 ;
        RECT 57.000 200.910 78.660 200.920 ;
        RECT 36.680 200.900 78.660 200.910 ;
        RECT 30.610 199.315 78.660 200.900 ;
        RECT 30.610 199.305 58.700 199.315 ;
        RECT 30.610 199.295 36.850 199.305 ;
        RECT 43.500 199.250 44.350 199.305 ;
        RECT 56.740 199.300 58.700 199.305 ;
        RECT 71.800 199.300 72.650 199.315 ;
      LAYER pwell ;
        RECT 36.550 199.015 37.000 199.100 ;
        RECT 39.400 199.015 40.100 199.050 ;
        RECT 30.815 199.000 33.545 199.005 ;
        RECT 30.815 198.905 34.000 199.000 ;
        RECT 36.550 198.915 40.100 199.015 ;
        RECT 42.650 199.015 44.150 199.100 ;
        RECT 46.700 199.015 47.350 199.100 ;
        RECT 42.650 198.915 47.350 199.015 ;
        RECT 49.850 199.015 50.750 199.100 ;
        RECT 53.300 199.015 53.900 199.150 ;
        RECT 49.850 198.915 53.900 199.015 ;
        RECT 56.450 199.025 58.300 199.100 ;
        RECT 60.750 199.025 61.500 199.150 ;
        RECT 56.450 198.925 61.500 199.025 ;
        RECT 64.000 199.025 64.850 199.150 ;
        RECT 67.400 199.025 68.100 199.100 ;
        RECT 64.000 198.925 68.100 199.025 ;
        RECT 70.600 199.025 72.450 199.100 ;
        RECT 75.000 199.025 75.800 199.050 ;
        RECT 70.600 198.925 75.800 199.025 ;
        RECT 56.450 198.915 78.465 198.925 ;
        RECT 36.550 198.905 78.465 198.915 ;
        RECT 30.815 198.200 78.465 198.905 ;
        RECT 30.815 198.150 64.145 198.200 ;
        RECT 30.815 198.105 39.615 198.150 ;
        RECT 40.005 198.105 42.755 198.150 ;
        RECT 44.105 198.105 46.835 198.150 ;
        RECT 47.255 198.105 50.005 198.150 ;
        RECT 50.655 198.105 53.385 198.150 ;
        RECT 53.805 198.105 56.555 198.150 ;
        RECT 58.205 198.115 60.935 198.150 ;
        RECT 61.395 198.115 64.145 198.150 ;
        RECT 64.755 198.150 78.465 198.200 ;
        RECT 64.755 198.115 67.485 198.150 ;
        RECT 67.945 198.115 70.695 198.150 ;
        RECT 72.365 198.115 75.095 198.150 ;
        RECT 75.715 198.115 78.465 198.150 ;
        RECT 30.815 198.100 37.000 198.105 ;
        RECT 30.815 198.095 33.545 198.100 ;
        RECT 33.905 198.095 36.655 198.100 ;
        RECT 30.945 197.905 31.115 198.095 ;
        RECT 34.045 197.905 34.215 198.095 ;
        RECT 37.015 197.915 37.185 198.105 ;
        RECT 40.145 197.915 40.315 198.105 ;
        RECT 44.235 197.915 44.405 198.105 ;
        RECT 47.395 197.915 47.565 198.105 ;
        RECT 50.785 197.915 50.955 198.105 ;
        RECT 53.945 197.915 54.115 198.105 ;
        RECT 58.335 197.925 58.505 198.115 ;
        RECT 61.535 197.925 61.705 198.115 ;
        RECT 64.885 197.925 65.055 198.115 ;
        RECT 68.085 197.925 68.255 198.115 ;
        RECT 72.495 197.925 72.665 198.115 ;
        RECT 75.855 197.925 76.025 198.115 ;
      LAYER nwell ;
        RECT 57.800 197.550 58.650 197.600 ;
        RECT 30.610 195.945 78.660 197.550 ;
        RECT 43.650 195.900 44.550 195.945 ;
        RECT 57.800 195.900 58.650 195.945 ;
      LAYER pwell ;
        RECT 33.900 195.655 34.550 195.700 ;
        RECT 40.000 195.655 40.750 195.700 ;
        RECT 47.200 195.655 47.700 195.700 ;
        RECT 53.750 195.655 54.350 195.700 ;
        RECT 61.300 195.655 62.000 195.700 ;
        RECT 67.850 195.655 68.500 195.700 ;
        RECT 30.845 195.555 34.550 195.655 ;
        RECT 36.915 195.555 40.750 195.655 ;
        RECT 44.135 195.650 47.700 195.655 ;
        RECT 42.400 195.555 47.700 195.650 ;
        RECT 50.685 195.600 54.350 195.655 ;
        RECT 58.235 195.650 62.000 195.655 ;
        RECT 50.250 195.555 54.350 195.600 ;
        RECT 56.900 195.555 62.000 195.650 ;
        RECT 64.785 195.600 68.500 195.655 ;
        RECT 64.550 195.555 68.500 195.600 ;
        RECT 71.050 195.655 72.500 195.700 ;
        RECT 75.450 195.655 76.750 195.700 ;
        RECT 71.050 195.555 76.750 195.655 ;
        RECT 30.845 195.500 36.275 195.555 ;
        RECT 36.915 195.500 78.465 195.555 ;
        RECT 30.845 194.850 78.465 195.500 ;
        RECT 30.845 194.745 34.015 194.850 ;
        RECT 34.445 194.745 36.275 194.850 ;
        RECT 36.915 194.800 56.995 194.850 ;
        RECT 57.205 194.830 57.635 194.850 ;
        RECT 36.915 194.745 40.085 194.800 ;
        RECT 40.665 194.745 42.495 194.800 ;
        RECT 44.135 194.745 47.305 194.800 ;
        RECT 47.605 194.745 50.355 194.800 ;
        RECT 50.685 194.745 53.855 194.800 ;
        RECT 54.245 194.745 56.995 194.800 ;
        RECT 58.235 194.800 64.645 194.850 ;
        RECT 58.235 194.745 61.405 194.800 ;
        RECT 61.895 194.745 64.645 194.800 ;
        RECT 64.785 194.800 78.465 194.850 ;
        RECT 64.785 194.745 67.955 194.800 ;
        RECT 68.395 194.745 71.145 194.800 ;
        RECT 72.385 194.745 75.555 194.800 ;
        RECT 76.635 194.745 78.465 194.800 ;
        RECT 30.945 194.555 31.115 194.745 ;
        RECT 34.585 194.555 34.755 194.745 ;
        RECT 37.015 194.555 37.185 194.745 ;
        RECT 40.805 194.555 40.975 194.745 ;
        RECT 44.235 194.555 44.405 194.745 ;
        RECT 47.745 194.555 47.915 194.745 ;
        RECT 50.785 194.555 50.955 194.745 ;
        RECT 54.385 194.555 54.555 194.745 ;
        RECT 58.335 194.555 58.505 194.745 ;
        RECT 62.035 194.555 62.205 194.745 ;
        RECT 64.885 194.555 65.055 194.745 ;
        RECT 68.535 194.555 68.705 194.745 ;
        RECT 72.485 194.555 72.655 194.745 ;
        RECT 76.775 194.555 76.945 194.745 ;
      LAYER li1 ;
        RECT 30.800 203.985 78.470 204.155 ;
        RECT 31.085 203.315 31.365 203.985 ;
        RECT 31.535 203.095 31.835 203.645 ;
        RECT 32.035 203.265 32.365 203.985 ;
        RECT 32.555 203.265 33.015 203.815 ;
        RECT 30.900 202.850 31.165 203.035 ;
        RECT 31.535 202.925 32.475 203.095 ;
        RECT 30.850 202.675 31.250 202.850 ;
        RECT 32.305 202.675 32.475 202.925 ;
        RECT 30.850 202.450 31.575 202.675 ;
        RECT 30.900 202.425 31.575 202.450 ;
        RECT 31.795 202.425 32.135 202.675 ;
        RECT 32.305 202.345 32.595 202.675 ;
        RECT 32.305 202.255 32.475 202.345 ;
        RECT 31.085 202.065 32.475 202.255 ;
        RECT 31.085 201.705 31.415 202.065 ;
        RECT 32.765 201.895 33.015 203.265 ;
        RECT 33.285 203.135 33.665 203.815 ;
        RECT 34.255 203.135 34.425 203.985 ;
        RECT 34.595 203.305 34.925 203.815 ;
        RECT 35.095 203.475 35.265 203.985 ;
        RECT 35.435 203.305 35.835 203.815 ;
        RECT 34.595 203.135 35.835 203.305 ;
        RECT 33.285 202.175 33.455 203.135 ;
        RECT 33.625 202.795 34.930 202.965 ;
        RECT 36.015 202.885 36.335 203.815 ;
        RECT 37.155 203.315 37.435 203.985 ;
        RECT 37.605 203.095 37.905 203.645 ;
        RECT 38.105 203.265 38.435 203.985 ;
        RECT 38.625 203.265 39.085 203.815 ;
        RECT 33.625 202.345 33.870 202.795 ;
        RECT 34.040 202.425 34.590 202.625 ;
        RECT 34.760 202.595 34.930 202.795 ;
        RECT 35.705 202.715 36.335 202.885 ;
        RECT 34.760 202.425 35.135 202.595 ;
        RECT 35.305 202.175 35.535 202.675 ;
        RECT 33.285 202.005 35.535 202.175 ;
        RECT 32.035 201.435 32.285 201.895 ;
        RECT 32.455 201.605 33.015 201.895 ;
        RECT 33.335 201.435 33.665 201.825 ;
        RECT 33.835 201.685 34.005 202.005 ;
        RECT 35.705 201.835 35.875 202.715 ;
        RECT 36.970 202.675 37.235 203.035 ;
        RECT 37.605 202.925 38.545 203.095 ;
        RECT 38.375 202.675 38.545 202.925 ;
        RECT 36.970 202.425 37.645 202.675 ;
        RECT 37.865 202.425 38.205 202.675 ;
        RECT 38.375 202.345 38.665 202.675 ;
        RECT 34.175 201.435 34.505 201.825 ;
        RECT 34.920 201.665 35.875 201.835 ;
        RECT 36.045 201.435 36.335 202.270 ;
        RECT 38.375 202.255 38.545 202.345 ;
        RECT 37.155 202.065 38.545 202.255 ;
        RECT 37.155 201.705 37.485 202.065 ;
        RECT 38.835 201.895 39.085 203.265 ;
        RECT 39.455 203.135 39.835 203.815 ;
        RECT 40.425 203.135 40.595 203.985 ;
        RECT 40.765 203.305 41.095 203.815 ;
        RECT 41.265 203.475 41.435 203.985 ;
        RECT 41.605 203.305 42.005 203.815 ;
        RECT 40.765 203.135 42.005 203.305 ;
        RECT 39.455 202.175 39.625 203.135 ;
        RECT 39.795 202.795 41.100 202.965 ;
        RECT 42.185 202.885 42.505 203.815 ;
        RECT 39.795 202.345 40.040 202.795 ;
        RECT 40.930 202.650 41.100 202.795 ;
        RECT 41.875 202.715 42.505 202.885 ;
        RECT 43.125 202.820 43.415 203.985 ;
        RECT 44.375 203.315 44.655 203.985 ;
        RECT 44.825 203.095 45.125 203.645 ;
        RECT 45.325 203.265 45.655 203.985 ;
        RECT 45.845 203.265 46.305 203.815 ;
        RECT 40.210 202.425 40.760 202.625 ;
        RECT 40.930 202.425 41.305 202.650 ;
        RECT 41.475 202.175 41.705 202.675 ;
        RECT 39.455 202.005 41.705 202.175 ;
        RECT 38.105 201.435 38.355 201.895 ;
        RECT 38.525 201.605 39.085 201.895 ;
        RECT 39.505 201.435 39.835 201.825 ;
        RECT 40.005 201.685 40.175 202.005 ;
        RECT 41.875 201.835 42.045 202.715 ;
        RECT 44.190 202.675 44.455 203.035 ;
        RECT 44.825 202.925 45.765 203.095 ;
        RECT 45.595 202.675 45.765 202.925 ;
        RECT 44.190 202.425 44.865 202.675 ;
        RECT 45.085 202.425 45.425 202.675 ;
        RECT 45.595 202.345 45.885 202.675 ;
        RECT 40.345 201.435 40.675 201.825 ;
        RECT 41.090 201.665 42.045 201.835 ;
        RECT 42.215 201.435 42.505 202.270 ;
        RECT 45.595 202.255 45.765 202.345 ;
        RECT 43.125 201.435 43.415 202.160 ;
        RECT 44.375 202.065 45.765 202.255 ;
        RECT 44.375 201.705 44.705 202.065 ;
        RECT 46.055 201.895 46.305 203.265 ;
        RECT 47.025 203.135 47.405 203.815 ;
        RECT 47.995 203.135 48.165 203.985 ;
        RECT 48.335 203.305 48.665 203.815 ;
        RECT 48.835 203.475 49.005 203.985 ;
        RECT 49.175 203.305 49.575 203.815 ;
        RECT 48.335 203.135 49.575 203.305 ;
        RECT 47.025 202.175 47.195 203.135 ;
        RECT 47.365 202.795 48.670 202.965 ;
        RECT 49.755 202.885 50.075 203.815 ;
        RECT 50.925 203.315 51.205 203.985 ;
        RECT 51.375 203.095 51.675 203.645 ;
        RECT 51.875 203.265 52.205 203.985 ;
        RECT 52.395 203.265 52.855 203.815 ;
        RECT 47.365 202.345 47.610 202.795 ;
        RECT 47.780 202.425 48.330 202.625 ;
        RECT 48.500 202.595 48.670 202.795 ;
        RECT 49.445 202.715 50.075 202.885 ;
        RECT 48.500 202.425 48.875 202.595 ;
        RECT 47.950 202.400 48.150 202.425 ;
        RECT 49.045 202.175 49.275 202.675 ;
        RECT 47.025 202.005 49.275 202.175 ;
        RECT 45.325 201.435 45.575 201.895 ;
        RECT 45.745 201.605 46.305 201.895 ;
        RECT 47.075 201.435 47.405 201.825 ;
        RECT 47.575 201.685 47.745 202.005 ;
        RECT 49.445 201.835 49.615 202.715 ;
        RECT 50.740 202.675 51.005 203.035 ;
        RECT 51.375 202.925 52.315 203.095 ;
        RECT 52.145 202.675 52.315 202.925 ;
        RECT 50.740 202.425 51.415 202.675 ;
        RECT 51.635 202.425 51.975 202.675 ;
        RECT 52.145 202.345 52.435 202.675 ;
        RECT 47.915 201.435 48.245 201.825 ;
        RECT 48.660 201.665 49.615 201.835 ;
        RECT 49.785 201.435 50.075 202.270 ;
        RECT 52.145 202.255 52.315 202.345 ;
        RECT 50.925 202.065 52.315 202.255 ;
        RECT 50.925 201.705 51.255 202.065 ;
        RECT 52.605 201.895 52.855 203.265 ;
        RECT 53.525 203.135 53.905 203.815 ;
        RECT 54.495 203.135 54.665 203.985 ;
        RECT 54.835 203.305 55.165 203.815 ;
        RECT 55.335 203.475 55.505 203.985 ;
        RECT 55.675 203.305 56.075 203.815 ;
        RECT 54.835 203.135 56.075 203.305 ;
        RECT 53.525 202.175 53.695 203.135 ;
        RECT 53.865 202.795 55.170 202.965 ;
        RECT 56.255 202.885 56.575 203.815 ;
        RECT 53.865 202.345 54.110 202.795 ;
        RECT 54.280 202.425 54.830 202.625 ;
        RECT 55.000 202.615 55.170 202.795 ;
        RECT 55.945 202.715 56.575 202.885 ;
        RECT 57.275 202.820 57.565 203.985 ;
        RECT 58.475 203.315 58.755 203.985 ;
        RECT 58.925 203.095 59.225 203.645 ;
        RECT 59.425 203.265 59.755 203.985 ;
        RECT 59.945 203.265 60.405 203.815 ;
        RECT 55.000 202.595 55.295 202.615 ;
        RECT 55.000 202.425 55.375 202.595 ;
        RECT 54.400 202.400 54.600 202.425 ;
        RECT 55.545 202.175 55.775 202.675 ;
        RECT 53.525 202.005 55.775 202.175 ;
        RECT 51.875 201.435 52.125 201.895 ;
        RECT 52.295 201.605 52.855 201.895 ;
        RECT 53.575 201.435 53.905 201.825 ;
        RECT 54.075 201.685 54.245 202.005 ;
        RECT 55.945 201.835 56.115 202.715 ;
        RECT 58.290 202.675 58.555 203.035 ;
        RECT 58.925 202.925 59.865 203.095 ;
        RECT 59.695 202.675 59.865 202.925 ;
        RECT 58.290 202.425 58.965 202.675 ;
        RECT 59.185 202.425 59.525 202.675 ;
        RECT 59.695 202.345 59.985 202.675 ;
        RECT 54.415 201.435 54.745 201.825 ;
        RECT 55.160 201.665 56.115 201.835 ;
        RECT 56.285 201.435 56.575 202.270 ;
        RECT 59.695 202.255 59.865 202.345 ;
        RECT 57.275 201.435 57.565 202.160 ;
        RECT 58.475 202.065 59.865 202.255 ;
        RECT 58.475 201.705 58.805 202.065 ;
        RECT 60.155 201.895 60.405 203.265 ;
        RECT 61.075 203.135 61.455 203.815 ;
        RECT 62.045 203.135 62.215 203.985 ;
        RECT 62.385 203.305 62.715 203.815 ;
        RECT 62.885 203.475 63.055 203.985 ;
        RECT 63.225 203.305 63.625 203.815 ;
        RECT 62.385 203.135 63.625 203.305 ;
        RECT 61.075 202.175 61.245 203.135 ;
        RECT 63.805 203.050 64.125 203.815 ;
        RECT 65.025 203.315 65.305 203.985 ;
        RECT 61.415 202.795 62.720 202.965 ;
        RECT 63.800 202.885 64.125 203.050 ;
        RECT 65.475 203.095 65.775 203.645 ;
        RECT 65.975 203.265 66.305 203.985 ;
        RECT 66.495 203.265 66.955 203.815 ;
        RECT 61.415 202.345 61.660 202.795 ;
        RECT 61.830 202.425 62.380 202.625 ;
        RECT 62.550 202.595 62.720 202.795 ;
        RECT 63.495 202.715 64.125 202.885 ;
        RECT 62.550 202.425 62.925 202.595 ;
        RECT 63.095 202.175 63.325 202.675 ;
        RECT 61.075 202.005 63.325 202.175 ;
        RECT 59.425 201.435 59.675 201.895 ;
        RECT 59.845 201.605 60.405 201.895 ;
        RECT 61.125 201.435 61.455 201.825 ;
        RECT 61.625 201.685 61.795 202.005 ;
        RECT 63.495 201.835 63.665 202.715 ;
        RECT 64.840 202.675 65.105 203.035 ;
        RECT 65.475 202.925 66.415 203.095 ;
        RECT 66.245 202.675 66.415 202.925 ;
        RECT 64.840 202.650 65.515 202.675 ;
        RECT 64.815 202.475 65.515 202.650 ;
        RECT 64.840 202.425 65.515 202.475 ;
        RECT 65.735 202.425 66.075 202.675 ;
        RECT 66.245 202.345 66.535 202.675 ;
        RECT 61.965 201.435 62.295 201.825 ;
        RECT 62.710 201.665 63.665 201.835 ;
        RECT 63.835 201.435 64.125 202.270 ;
        RECT 66.245 202.255 66.415 202.345 ;
        RECT 65.025 202.065 66.415 202.255 ;
        RECT 65.025 201.705 65.355 202.065 ;
        RECT 66.705 201.895 66.955 203.265 ;
        RECT 67.625 203.135 68.005 203.815 ;
        RECT 68.595 203.135 68.765 203.985 ;
        RECT 68.935 203.305 69.265 203.815 ;
        RECT 69.435 203.475 69.605 203.985 ;
        RECT 69.775 203.305 70.175 203.815 ;
        RECT 68.935 203.135 70.175 203.305 ;
        RECT 67.625 202.175 67.795 203.135 ;
        RECT 67.965 202.795 69.270 202.965 ;
        RECT 70.355 202.885 70.675 203.815 ;
        RECT 67.965 202.345 68.210 202.795 ;
        RECT 68.380 202.425 68.930 202.625 ;
        RECT 69.100 202.595 69.270 202.795 ;
        RECT 70.045 202.715 70.675 202.885 ;
        RECT 71.385 202.820 71.675 203.985 ;
        RECT 72.635 203.315 72.915 203.985 ;
        RECT 73.085 203.095 73.385 203.645 ;
        RECT 73.585 203.265 73.915 203.985 ;
        RECT 74.105 203.265 74.565 203.815 ;
        RECT 69.100 202.425 69.475 202.595 ;
        RECT 69.645 202.175 69.875 202.675 ;
        RECT 67.625 202.005 69.875 202.175 ;
        RECT 65.975 201.435 66.225 201.895 ;
        RECT 66.395 201.605 66.955 201.895 ;
        RECT 67.675 201.435 68.005 201.825 ;
        RECT 68.175 201.685 68.345 202.005 ;
        RECT 70.045 201.835 70.215 202.715 ;
        RECT 72.450 202.675 72.715 203.035 ;
        RECT 73.085 202.925 74.025 203.095 ;
        RECT 73.855 202.675 74.025 202.925 ;
        RECT 72.450 202.425 73.125 202.675 ;
        RECT 73.345 202.425 73.685 202.675 ;
        RECT 73.855 202.345 74.145 202.675 ;
        RECT 68.515 201.435 68.845 201.825 ;
        RECT 69.260 201.665 70.215 201.835 ;
        RECT 70.385 201.435 70.675 202.270 ;
        RECT 73.855 202.255 74.025 202.345 ;
        RECT 71.385 201.435 71.675 202.160 ;
        RECT 72.635 202.065 74.025 202.255 ;
        RECT 72.635 201.705 72.965 202.065 ;
        RECT 74.315 201.895 74.565 203.265 ;
        RECT 75.335 203.135 75.715 203.815 ;
        RECT 76.305 203.135 76.475 203.985 ;
        RECT 76.645 203.305 76.975 203.815 ;
        RECT 77.145 203.475 77.315 203.985 ;
        RECT 77.485 203.305 77.885 203.815 ;
        RECT 76.645 203.135 77.885 203.305 ;
        RECT 75.335 202.175 75.505 203.135 ;
        RECT 75.675 202.795 76.980 202.965 ;
        RECT 78.065 202.885 78.385 203.815 ;
        RECT 75.675 202.345 75.920 202.795 ;
        RECT 76.090 202.425 76.640 202.625 ;
        RECT 76.810 202.600 76.980 202.795 ;
        RECT 77.755 202.715 78.385 202.885 ;
        RECT 76.810 202.595 77.100 202.600 ;
        RECT 76.810 202.425 77.185 202.595 ;
        RECT 76.900 202.400 77.100 202.425 ;
        RECT 77.355 202.175 77.585 202.675 ;
        RECT 75.335 202.005 77.585 202.175 ;
        RECT 73.585 201.435 73.835 201.895 ;
        RECT 74.005 201.605 74.565 201.895 ;
        RECT 75.385 201.435 75.715 201.825 ;
        RECT 75.885 201.685 76.055 202.005 ;
        RECT 77.755 201.835 77.925 202.715 ;
        RECT 76.225 201.435 76.555 201.825 ;
        RECT 76.970 201.665 77.925 201.835 ;
        RECT 78.095 201.435 78.385 202.270 ;
        RECT 30.800 201.265 78.470 201.435 ;
        RECT 39.080 201.260 39.400 201.265 ;
        RECT 56.350 200.815 57.200 200.830 ;
        RECT 56.350 200.805 78.470 200.815 ;
        RECT 36.645 200.795 78.470 200.805 ;
        RECT 30.800 200.645 78.470 200.795 ;
        RECT 30.800 200.635 56.560 200.645 ;
        RECT 30.800 200.625 36.955 200.635 ;
        RECT 30.895 198.255 31.155 200.445 ;
        RECT 31.325 199.895 31.665 200.625 ;
        RECT 31.845 199.715 32.115 200.445 ;
        RECT 31.345 199.495 32.115 199.715 ;
        RECT 32.295 199.735 32.525 200.445 ;
        RECT 32.695 199.915 33.025 200.625 ;
        RECT 33.195 199.735 33.455 200.445 ;
        RECT 32.295 199.495 33.455 199.735 ;
        RECT 33.985 199.535 36.575 200.625 ;
        RECT 31.345 198.825 31.635 199.495 ;
        RECT 31.815 199.005 32.280 199.315 ;
        RECT 32.460 199.005 32.985 199.315 ;
        RECT 31.345 198.625 32.575 198.825 ;
        RECT 32.755 198.700 32.985 199.005 ;
        RECT 33.165 198.985 33.465 199.315 ;
        RECT 33.985 198.845 35.195 199.365 ;
        RECT 35.365 199.015 36.575 199.535 ;
        RECT 31.415 198.075 32.085 198.445 ;
        RECT 32.265 198.255 32.575 198.625 ;
        RECT 32.750 198.500 32.985 198.700 ;
        RECT 32.755 198.365 32.985 198.500 ;
        RECT 33.165 198.075 33.455 198.805 ;
        RECT 33.985 198.100 36.575 198.845 ;
        RECT 36.965 198.265 37.225 200.455 ;
        RECT 37.395 199.905 37.735 200.635 ;
        RECT 37.915 199.725 38.185 200.455 ;
        RECT 37.415 199.505 38.185 199.725 ;
        RECT 38.365 199.745 38.595 200.455 ;
        RECT 38.765 199.925 39.095 200.635 ;
        RECT 39.265 199.745 39.525 200.455 ;
        RECT 38.365 199.505 39.525 199.745 ;
        RECT 40.085 199.545 42.675 200.635 ;
        RECT 37.415 198.835 37.705 199.505 ;
        RECT 37.885 199.015 38.350 199.325 ;
        RECT 38.530 199.015 39.055 199.325 ;
        RECT 37.415 198.635 38.645 198.835 ;
        RECT 33.985 198.085 36.900 198.100 ;
        RECT 37.485 198.085 38.155 198.455 ;
        RECT 38.335 198.265 38.645 198.635 ;
        RECT 38.825 198.375 39.055 199.015 ;
        RECT 39.235 198.995 39.535 199.325 ;
        RECT 40.085 198.855 41.295 199.375 ;
        RECT 41.465 199.025 42.675 199.545 ;
        RECT 43.125 199.470 43.415 200.635 ;
        RECT 39.235 198.085 39.525 198.815 ;
        RECT 40.085 198.085 42.675 198.855 ;
        RECT 43.125 198.085 43.415 198.810 ;
        RECT 44.185 198.265 44.445 200.455 ;
        RECT 44.615 199.905 44.955 200.635 ;
        RECT 45.135 199.725 45.405 200.455 ;
        RECT 44.635 199.505 45.405 199.725 ;
        RECT 45.585 199.745 45.815 200.455 ;
        RECT 45.985 199.925 46.315 200.635 ;
        RECT 46.485 199.745 46.745 200.455 ;
        RECT 45.585 199.505 46.745 199.745 ;
        RECT 47.335 199.545 49.925 200.635 ;
        RECT 44.635 198.835 44.925 199.505 ;
        RECT 45.105 199.015 45.570 199.325 ;
        RECT 45.750 199.015 46.275 199.325 ;
        RECT 44.635 198.635 45.865 198.835 ;
        RECT 44.705 198.085 45.375 198.455 ;
        RECT 45.555 198.265 45.865 198.635 ;
        RECT 46.045 198.375 46.275 199.015 ;
        RECT 46.455 198.995 46.755 199.325 ;
        RECT 47.335 198.855 48.545 199.375 ;
        RECT 48.715 199.025 49.925 199.545 ;
        RECT 46.455 198.085 46.745 198.815 ;
        RECT 47.335 198.085 49.925 198.855 ;
        RECT 50.735 198.265 50.995 200.455 ;
        RECT 51.165 199.905 51.505 200.635 ;
        RECT 51.685 199.725 51.955 200.455 ;
        RECT 51.185 199.505 51.955 199.725 ;
        RECT 52.135 199.745 52.365 200.455 ;
        RECT 52.535 199.925 52.865 200.635 ;
        RECT 53.035 199.745 53.295 200.455 ;
        RECT 52.135 199.505 53.295 199.745 ;
        RECT 53.885 199.545 56.475 200.635 ;
        RECT 51.185 198.835 51.475 199.505 ;
        RECT 51.655 199.015 52.120 199.325 ;
        RECT 52.300 199.015 52.825 199.325 ;
        RECT 51.185 198.635 52.415 198.835 ;
        RECT 51.255 198.085 51.925 198.455 ;
        RECT 52.105 198.265 52.415 198.635 ;
        RECT 52.595 198.375 52.825 199.015 ;
        RECT 53.005 198.995 53.305 199.325 ;
        RECT 53.885 198.855 55.095 199.375 ;
        RECT 55.265 199.025 56.475 199.545 ;
        RECT 57.275 199.480 57.565 200.645 ;
        RECT 53.005 198.085 53.295 198.815 ;
        RECT 53.885 198.095 56.475 198.855 ;
        RECT 57.275 198.095 57.565 198.820 ;
        RECT 58.285 198.275 58.545 200.465 ;
        RECT 58.715 199.915 59.055 200.645 ;
        RECT 59.235 199.735 59.505 200.465 ;
        RECT 58.735 199.515 59.505 199.735 ;
        RECT 59.685 199.755 59.915 200.465 ;
        RECT 60.085 199.935 60.415 200.645 ;
        RECT 60.585 199.755 60.845 200.465 ;
        RECT 59.685 199.515 60.845 199.755 ;
        RECT 61.475 199.555 64.065 200.645 ;
        RECT 58.735 198.845 59.025 199.515 ;
        RECT 59.205 199.025 59.670 199.335 ;
        RECT 59.850 199.025 60.375 199.335 ;
        RECT 58.735 198.645 59.965 198.845 ;
        RECT 58.805 198.095 59.475 198.465 ;
        RECT 59.655 198.275 59.965 198.645 ;
        RECT 60.145 198.385 60.375 199.025 ;
        RECT 60.555 199.005 60.855 199.335 ;
        RECT 61.475 198.865 62.685 199.385 ;
        RECT 62.855 199.035 64.065 199.555 ;
        RECT 60.555 198.095 60.845 198.825 ;
        RECT 61.475 198.095 64.065 198.865 ;
        RECT 64.835 198.275 65.095 200.465 ;
        RECT 65.265 199.915 65.605 200.645 ;
        RECT 65.785 199.735 66.055 200.465 ;
        RECT 65.285 199.515 66.055 199.735 ;
        RECT 66.235 199.755 66.465 200.465 ;
        RECT 66.635 199.935 66.965 200.645 ;
        RECT 67.135 199.755 67.395 200.465 ;
        RECT 66.235 199.515 67.395 199.755 ;
        RECT 68.025 199.555 70.615 200.645 ;
        RECT 65.285 198.845 65.575 199.515 ;
        RECT 65.755 199.025 66.220 199.335 ;
        RECT 66.400 199.025 66.925 199.335 ;
        RECT 65.285 198.645 66.515 198.845 ;
        RECT 65.355 198.095 66.025 198.465 ;
        RECT 66.205 198.275 66.515 198.645 ;
        RECT 66.695 198.385 66.925 199.025 ;
        RECT 67.105 199.005 67.405 199.335 ;
        RECT 68.025 198.865 69.235 199.385 ;
        RECT 69.405 199.035 70.615 199.555 ;
        RECT 71.385 199.480 71.675 200.645 ;
        RECT 67.105 198.095 67.395 198.825 ;
        RECT 68.025 198.095 70.615 198.865 ;
        RECT 71.385 198.095 71.675 198.820 ;
        RECT 72.445 198.275 72.705 200.465 ;
        RECT 72.875 199.915 73.215 200.645 ;
        RECT 73.395 199.735 73.665 200.465 ;
        RECT 72.895 199.515 73.665 199.735 ;
        RECT 73.845 199.755 74.075 200.465 ;
        RECT 74.245 199.935 74.575 200.645 ;
        RECT 74.745 199.755 75.005 200.465 ;
        RECT 73.845 199.515 75.005 199.755 ;
        RECT 75.795 199.555 78.385 200.645 ;
        RECT 72.895 198.845 73.185 199.515 ;
        RECT 73.365 199.025 73.830 199.335 ;
        RECT 74.010 199.025 74.535 199.335 ;
        RECT 72.895 198.645 74.125 198.845 ;
        RECT 72.965 198.095 73.635 198.465 ;
        RECT 73.815 198.275 74.125 198.645 ;
        RECT 74.305 198.385 74.535 199.025 ;
        RECT 74.715 199.005 75.015 199.335 ;
        RECT 75.795 198.865 77.005 199.385 ;
        RECT 77.175 199.035 78.385 199.555 ;
        RECT 74.715 198.095 75.005 198.825 ;
        RECT 75.795 198.095 78.385 198.865 ;
        RECT 53.885 198.085 78.470 198.095 ;
        RECT 33.985 198.075 78.470 198.085 ;
        RECT 30.800 197.925 78.470 198.075 ;
        RECT 30.800 197.920 57.225 197.925 ;
        RECT 60.935 197.920 61.430 197.925 ;
        RECT 30.800 197.915 57.205 197.920 ;
        RECT 30.800 197.905 36.660 197.915 ;
        RECT 30.800 197.275 78.470 197.445 ;
        RECT 30.885 196.425 31.265 197.105 ;
        RECT 31.855 196.425 32.025 197.275 ;
        RECT 32.195 196.595 32.525 197.105 ;
        RECT 32.695 196.765 32.865 197.275 ;
        RECT 33.035 196.595 33.435 197.105 ;
        RECT 32.195 196.425 33.435 196.595 ;
        RECT 30.885 195.465 31.055 196.425 ;
        RECT 31.225 196.085 32.530 196.255 ;
        RECT 33.615 196.175 33.935 197.105 ;
        RECT 34.525 196.185 36.195 197.275 ;
        RECT 31.225 195.635 31.470 196.085 ;
        RECT 31.640 195.715 32.190 195.915 ;
        RECT 32.360 195.885 32.530 196.085 ;
        RECT 33.305 196.005 33.935 196.175 ;
        RECT 32.360 195.715 32.735 195.885 ;
        RECT 32.905 195.465 33.135 195.965 ;
        RECT 30.885 195.295 33.135 195.465 ;
        RECT 30.935 194.725 31.265 195.115 ;
        RECT 31.435 194.975 31.605 195.295 ;
        RECT 33.305 195.125 33.475 196.005 ;
        RECT 31.775 194.725 32.105 195.115 ;
        RECT 32.520 194.955 33.475 195.125 ;
        RECT 33.645 194.725 33.935 195.560 ;
        RECT 34.525 195.495 35.275 196.015 ;
        RECT 35.445 195.665 36.195 196.185 ;
        RECT 36.955 196.425 37.335 197.105 ;
        RECT 37.925 196.425 38.095 197.275 ;
        RECT 38.265 196.595 38.595 197.105 ;
        RECT 38.765 196.765 38.935 197.275 ;
        RECT 39.105 196.595 39.505 197.105 ;
        RECT 38.265 196.425 39.505 196.595 ;
        RECT 34.525 194.725 36.195 195.495 ;
        RECT 36.955 195.465 37.125 196.425 ;
        RECT 37.295 196.085 38.600 196.255 ;
        RECT 39.685 196.175 40.005 197.105 ;
        RECT 40.745 196.185 42.415 197.275 ;
        RECT 37.295 195.635 37.540 196.085 ;
        RECT 37.710 195.715 38.260 195.915 ;
        RECT 38.430 195.885 38.600 196.085 ;
        RECT 39.375 196.005 40.005 196.175 ;
        RECT 38.430 195.715 38.805 195.885 ;
        RECT 38.975 195.465 39.205 195.965 ;
        RECT 36.955 195.295 39.205 195.465 ;
        RECT 37.005 194.725 37.335 195.115 ;
        RECT 37.505 194.975 37.675 195.295 ;
        RECT 39.375 195.125 39.545 196.005 ;
        RECT 37.845 194.725 38.175 195.115 ;
        RECT 38.590 194.955 39.545 195.125 ;
        RECT 39.715 194.725 40.005 195.560 ;
        RECT 40.745 195.495 41.495 196.015 ;
        RECT 41.665 195.665 42.415 196.185 ;
        RECT 43.125 196.110 43.415 197.275 ;
        RECT 44.175 196.425 44.555 197.105 ;
        RECT 45.145 196.425 45.315 197.275 ;
        RECT 45.485 196.595 45.815 197.105 ;
        RECT 45.985 196.765 46.155 197.275 ;
        RECT 46.325 196.595 46.725 197.105 ;
        RECT 45.485 196.425 46.725 196.595 ;
        RECT 40.745 194.725 42.415 195.495 ;
        RECT 44.175 195.465 44.345 196.425 ;
        RECT 44.515 196.085 45.820 196.255 ;
        RECT 46.905 196.175 47.225 197.105 ;
        RECT 47.685 196.185 50.275 197.275 ;
        RECT 44.515 195.635 44.760 196.085 ;
        RECT 44.930 195.715 45.480 195.915 ;
        RECT 45.650 195.885 45.820 196.085 ;
        RECT 46.595 196.005 47.225 196.175 ;
        RECT 45.650 195.715 46.025 195.885 ;
        RECT 46.195 195.465 46.425 195.965 ;
        RECT 43.125 194.725 43.415 195.450 ;
        RECT 44.175 195.295 46.425 195.465 ;
        RECT 44.225 194.725 44.555 195.115 ;
        RECT 44.725 194.975 44.895 195.295 ;
        RECT 46.595 195.125 46.765 196.005 ;
        RECT 45.065 194.725 45.395 195.115 ;
        RECT 45.810 194.955 46.765 195.125 ;
        RECT 46.935 194.725 47.225 195.560 ;
        RECT 47.685 195.495 48.895 196.015 ;
        RECT 49.065 195.665 50.275 196.185 ;
        RECT 50.725 196.425 51.105 197.105 ;
        RECT 51.695 196.425 51.865 197.275 ;
        RECT 52.035 196.595 52.365 197.105 ;
        RECT 52.535 196.765 52.705 197.275 ;
        RECT 52.875 196.595 53.275 197.105 ;
        RECT 52.035 196.425 53.275 196.595 ;
        RECT 47.685 194.725 50.275 195.495 ;
        RECT 50.725 195.465 50.895 196.425 ;
        RECT 51.065 196.085 52.370 196.255 ;
        RECT 53.455 196.175 53.775 197.105 ;
        RECT 54.325 196.185 56.915 197.275 ;
        RECT 51.065 195.635 51.310 196.085 ;
        RECT 51.480 195.715 52.030 195.915 ;
        RECT 52.200 195.885 52.370 196.085 ;
        RECT 53.145 196.005 53.775 196.175 ;
        RECT 52.200 195.715 52.575 195.885 ;
        RECT 52.745 195.465 52.975 195.965 ;
        RECT 50.725 195.295 52.975 195.465 ;
        RECT 50.775 194.725 51.105 195.115 ;
        RECT 51.275 194.975 51.445 195.295 ;
        RECT 53.145 195.125 53.315 196.005 ;
        RECT 51.615 194.725 51.945 195.115 ;
        RECT 52.360 194.955 53.315 195.125 ;
        RECT 53.485 194.725 53.775 195.560 ;
        RECT 54.325 195.495 55.535 196.015 ;
        RECT 55.705 195.665 56.915 196.185 ;
        RECT 57.275 196.110 57.565 197.275 ;
        RECT 58.275 196.425 58.655 197.105 ;
        RECT 59.245 196.425 59.415 197.275 ;
        RECT 59.585 196.595 59.915 197.105 ;
        RECT 60.085 196.765 60.255 197.275 ;
        RECT 60.425 196.595 60.825 197.105 ;
        RECT 59.585 196.425 60.825 196.595 ;
        RECT 54.325 194.725 56.915 195.495 ;
        RECT 58.275 195.465 58.445 196.425 ;
        RECT 58.615 196.085 59.920 196.255 ;
        RECT 61.005 196.175 61.325 197.105 ;
        RECT 61.975 196.185 64.565 197.275 ;
        RECT 58.615 195.635 58.860 196.085 ;
        RECT 59.030 195.715 59.580 195.915 ;
        RECT 59.750 195.885 59.920 196.085 ;
        RECT 60.695 196.005 61.325 196.175 ;
        RECT 59.750 195.715 60.125 195.885 ;
        RECT 60.295 195.465 60.525 195.965 ;
        RECT 57.275 194.725 57.565 195.450 ;
        RECT 58.275 195.295 60.525 195.465 ;
        RECT 58.325 194.725 58.655 195.115 ;
        RECT 58.825 194.975 58.995 195.295 ;
        RECT 60.695 195.125 60.865 196.005 ;
        RECT 59.165 194.725 59.495 195.115 ;
        RECT 59.910 194.955 60.865 195.125 ;
        RECT 61.035 194.725 61.325 195.560 ;
        RECT 61.975 195.495 63.185 196.015 ;
        RECT 63.355 195.665 64.565 196.185 ;
        RECT 64.825 196.425 65.205 197.105 ;
        RECT 65.795 196.425 65.965 197.275 ;
        RECT 66.135 196.595 66.465 197.105 ;
        RECT 66.635 196.765 66.805 197.275 ;
        RECT 66.975 196.595 67.375 197.105 ;
        RECT 66.135 196.425 67.375 196.595 ;
        RECT 61.975 194.725 64.565 195.495 ;
        RECT 64.825 195.465 64.995 196.425 ;
        RECT 65.165 196.085 66.470 196.255 ;
        RECT 67.555 196.175 67.875 197.105 ;
        RECT 68.475 196.185 71.065 197.275 ;
        RECT 65.165 195.635 65.410 196.085 ;
        RECT 65.580 195.715 66.130 195.915 ;
        RECT 66.300 195.885 66.470 196.085 ;
        RECT 67.245 196.005 67.875 196.175 ;
        RECT 66.300 195.715 66.675 195.885 ;
        RECT 66.845 195.465 67.075 195.965 ;
        RECT 64.825 195.295 67.075 195.465 ;
        RECT 64.875 194.725 65.205 195.115 ;
        RECT 65.375 194.975 65.545 195.295 ;
        RECT 67.245 195.125 67.415 196.005 ;
        RECT 65.715 194.725 66.045 195.115 ;
        RECT 66.460 194.955 67.415 195.125 ;
        RECT 67.585 194.725 67.875 195.560 ;
        RECT 68.475 195.495 69.685 196.015 ;
        RECT 69.855 195.665 71.065 196.185 ;
        RECT 71.385 196.110 71.675 197.275 ;
        RECT 72.425 196.425 72.805 197.105 ;
        RECT 73.395 196.425 73.565 197.275 ;
        RECT 73.735 196.595 74.065 197.105 ;
        RECT 74.235 196.765 74.405 197.275 ;
        RECT 74.575 196.595 74.975 197.105 ;
        RECT 73.735 196.425 74.975 196.595 ;
        RECT 68.475 194.725 71.065 195.495 ;
        RECT 72.425 195.465 72.595 196.425 ;
        RECT 72.765 196.085 74.070 196.255 ;
        RECT 75.155 196.175 75.475 197.105 ;
        RECT 76.715 196.185 78.385 197.275 ;
        RECT 72.765 195.635 73.010 196.085 ;
        RECT 73.180 195.715 73.730 195.915 ;
        RECT 73.900 195.885 74.070 196.085 ;
        RECT 74.845 196.005 75.475 196.175 ;
        RECT 73.900 195.715 74.275 195.885 ;
        RECT 74.445 195.465 74.675 195.965 ;
        RECT 71.385 194.725 71.675 195.450 ;
        RECT 72.425 195.295 74.675 195.465 ;
        RECT 72.475 194.725 72.805 195.115 ;
        RECT 72.975 194.975 73.145 195.295 ;
        RECT 74.845 195.125 75.015 196.005 ;
        RECT 73.315 194.725 73.645 195.115 ;
        RECT 74.060 194.955 75.015 195.125 ;
        RECT 75.185 194.725 75.475 195.560 ;
        RECT 76.715 195.495 77.465 196.015 ;
        RECT 77.635 195.665 78.385 196.185 ;
        RECT 76.715 194.725 78.385 195.495 ;
        RECT 30.800 194.555 78.470 194.725 ;
        RECT 50.310 194.550 50.670 194.555 ;
      LAYER mcon ;
        RECT 30.945 203.985 31.115 204.155 ;
        RECT 31.405 203.985 31.575 204.155 ;
        RECT 31.865 203.985 32.035 204.155 ;
        RECT 32.325 203.985 32.495 204.155 ;
        RECT 32.785 203.985 32.955 204.155 ;
        RECT 33.345 203.985 33.515 204.155 ;
        RECT 33.805 203.985 33.975 204.155 ;
        RECT 34.265 203.985 34.435 204.155 ;
        RECT 34.725 203.985 34.895 204.155 ;
        RECT 35.185 203.985 35.355 204.155 ;
        RECT 35.645 203.985 35.815 204.155 ;
        RECT 36.105 203.985 36.275 204.155 ;
        RECT 37.015 203.985 37.185 204.155 ;
        RECT 37.475 203.985 37.645 204.155 ;
        RECT 37.935 203.985 38.105 204.155 ;
        RECT 38.395 203.985 38.565 204.155 ;
        RECT 38.855 203.985 39.025 204.155 ;
        RECT 39.515 203.985 39.685 204.155 ;
        RECT 39.975 203.985 40.145 204.155 ;
        RECT 40.435 203.985 40.605 204.155 ;
        RECT 40.895 203.985 41.065 204.155 ;
        RECT 41.355 203.985 41.525 204.155 ;
        RECT 41.815 203.985 41.985 204.155 ;
        RECT 42.275 203.985 42.445 204.155 ;
        RECT 43.185 203.985 43.355 204.155 ;
        RECT 44.235 203.985 44.405 204.155 ;
        RECT 44.695 203.985 44.865 204.155 ;
        RECT 45.155 203.985 45.325 204.155 ;
        RECT 45.615 203.985 45.785 204.155 ;
        RECT 46.075 203.985 46.245 204.155 ;
        RECT 47.085 203.985 47.255 204.155 ;
        RECT 47.545 203.985 47.715 204.155 ;
        RECT 48.005 203.985 48.175 204.155 ;
        RECT 48.465 203.985 48.635 204.155 ;
        RECT 48.925 203.985 49.095 204.155 ;
        RECT 49.385 203.985 49.555 204.155 ;
        RECT 49.845 203.985 50.015 204.155 ;
        RECT 50.785 203.985 50.955 204.155 ;
        RECT 51.245 203.985 51.415 204.155 ;
        RECT 51.705 203.985 51.875 204.155 ;
        RECT 52.165 203.985 52.335 204.155 ;
        RECT 52.625 203.985 52.795 204.155 ;
        RECT 53.585 203.985 53.755 204.155 ;
        RECT 54.045 203.985 54.215 204.155 ;
        RECT 54.505 203.985 54.675 204.155 ;
        RECT 54.965 203.985 55.135 204.155 ;
        RECT 55.425 203.985 55.595 204.155 ;
        RECT 55.885 203.985 56.055 204.155 ;
        RECT 56.345 203.985 56.515 204.155 ;
        RECT 57.335 203.985 57.505 204.155 ;
        RECT 58.335 203.985 58.505 204.155 ;
        RECT 58.795 203.985 58.965 204.155 ;
        RECT 59.255 203.985 59.425 204.155 ;
        RECT 59.715 203.985 59.885 204.155 ;
        RECT 60.175 203.985 60.345 204.155 ;
        RECT 61.135 203.985 61.305 204.155 ;
        RECT 61.595 203.985 61.765 204.155 ;
        RECT 62.055 203.985 62.225 204.155 ;
        RECT 62.515 203.985 62.685 204.155 ;
        RECT 62.975 203.985 63.145 204.155 ;
        RECT 63.435 203.985 63.605 204.155 ;
        RECT 63.895 203.985 64.065 204.155 ;
        RECT 64.885 203.985 65.055 204.155 ;
        RECT 65.345 203.985 65.515 204.155 ;
        RECT 65.805 203.985 65.975 204.155 ;
        RECT 66.265 203.985 66.435 204.155 ;
        RECT 66.725 203.985 66.895 204.155 ;
        RECT 67.685 203.985 67.855 204.155 ;
        RECT 68.145 203.985 68.315 204.155 ;
        RECT 68.605 203.985 68.775 204.155 ;
        RECT 69.065 203.985 69.235 204.155 ;
        RECT 69.525 203.985 69.695 204.155 ;
        RECT 69.985 203.985 70.155 204.155 ;
        RECT 70.445 203.985 70.615 204.155 ;
        RECT 71.445 203.985 71.615 204.155 ;
        RECT 72.495 203.985 72.665 204.155 ;
        RECT 72.955 203.985 73.125 204.155 ;
        RECT 73.415 203.985 73.585 204.155 ;
        RECT 73.875 203.985 74.045 204.155 ;
        RECT 74.335 203.985 74.505 204.155 ;
        RECT 75.395 203.985 75.565 204.155 ;
        RECT 75.855 203.985 76.025 204.155 ;
        RECT 76.315 203.985 76.485 204.155 ;
        RECT 76.775 203.985 76.945 204.155 ;
        RECT 77.235 203.985 77.405 204.155 ;
        RECT 77.695 203.985 77.865 204.155 ;
        RECT 78.155 203.985 78.325 204.155 ;
        RECT 30.950 202.550 31.150 202.750 ;
        RECT 31.850 202.450 32.050 202.650 ;
        RECT 32.785 202.115 32.955 202.285 ;
        RECT 33.655 202.700 33.830 202.880 ;
        RECT 34.200 202.440 34.380 202.615 ;
        RECT 36.105 202.795 36.275 202.965 ;
        RECT 37.000 202.500 37.200 202.700 ;
        RECT 37.945 202.425 38.115 202.595 ;
        RECT 38.850 202.050 39.050 202.250 ;
        RECT 42.275 202.795 42.445 202.965 ;
        RECT 40.375 202.425 40.550 202.605 ;
        RECT 41.055 202.425 41.225 202.595 ;
        RECT 44.250 202.450 44.450 202.650 ;
        RECT 45.165 202.465 45.335 202.640 ;
        RECT 46.085 202.455 46.260 202.625 ;
        RECT 47.400 202.425 47.580 202.600 ;
        RECT 49.850 202.800 50.050 203.000 ;
        RECT 50.750 202.450 50.950 202.650 ;
        RECT 51.705 202.455 51.875 202.625 ;
        RECT 52.650 202.350 52.820 202.520 ;
        RECT 56.275 202.885 56.445 203.055 ;
        RECT 55.125 202.440 55.295 202.615 ;
        RECT 58.335 202.465 58.505 202.640 ;
        RECT 59.250 202.450 59.450 202.650 ;
        RECT 60.200 202.650 60.370 202.825 ;
        RECT 62.000 202.425 62.170 202.595 ;
        RECT 63.800 202.850 64.000 203.050 ;
        RECT 62.675 202.425 62.845 202.595 ;
        RECT 65.805 202.455 65.975 202.625 ;
        RECT 66.725 202.395 66.895 202.575 ;
        RECT 67.965 202.425 68.135 202.595 ;
        RECT 68.550 202.435 68.720 202.610 ;
        RECT 70.400 202.800 70.600 203.000 ;
        RECT 74.200 203.300 74.400 203.500 ;
        RECT 72.495 202.455 72.665 202.625 ;
        RECT 73.425 202.425 73.595 202.595 ;
        RECT 76.260 202.425 76.430 202.595 ;
        RECT 78.100 202.800 78.300 203.000 ;
        RECT 30.945 201.265 31.115 201.435 ;
        RECT 31.405 201.265 31.575 201.435 ;
        RECT 31.865 201.265 32.035 201.435 ;
        RECT 32.325 201.265 32.495 201.435 ;
        RECT 32.785 201.265 32.955 201.435 ;
        RECT 33.345 201.265 33.515 201.435 ;
        RECT 33.805 201.265 33.975 201.435 ;
        RECT 34.265 201.265 34.435 201.435 ;
        RECT 34.725 201.265 34.895 201.435 ;
        RECT 35.185 201.265 35.355 201.435 ;
        RECT 35.645 201.265 35.815 201.435 ;
        RECT 36.105 201.265 36.275 201.435 ;
        RECT 37.015 201.265 37.185 201.435 ;
        RECT 37.475 201.265 37.645 201.435 ;
        RECT 37.935 201.265 38.105 201.435 ;
        RECT 38.395 201.265 38.565 201.435 ;
        RECT 38.855 201.265 39.025 201.435 ;
        RECT 39.515 201.265 39.685 201.435 ;
        RECT 39.975 201.265 40.145 201.435 ;
        RECT 40.435 201.265 40.605 201.435 ;
        RECT 40.895 201.265 41.065 201.435 ;
        RECT 41.355 201.265 41.525 201.435 ;
        RECT 41.815 201.265 41.985 201.435 ;
        RECT 42.275 201.265 42.445 201.435 ;
        RECT 43.185 201.265 43.355 201.435 ;
        RECT 44.235 201.265 44.405 201.435 ;
        RECT 44.695 201.265 44.865 201.435 ;
        RECT 45.155 201.265 45.325 201.435 ;
        RECT 45.615 201.265 45.785 201.435 ;
        RECT 46.075 201.265 46.245 201.435 ;
        RECT 47.085 201.265 47.255 201.435 ;
        RECT 47.545 201.265 47.715 201.435 ;
        RECT 48.005 201.265 48.175 201.435 ;
        RECT 48.465 201.265 48.635 201.435 ;
        RECT 48.925 201.265 49.095 201.435 ;
        RECT 49.385 201.265 49.555 201.435 ;
        RECT 49.845 201.265 50.015 201.435 ;
        RECT 50.785 201.265 50.955 201.435 ;
        RECT 51.245 201.265 51.415 201.435 ;
        RECT 51.705 201.265 51.875 201.435 ;
        RECT 52.165 201.265 52.335 201.435 ;
        RECT 52.625 201.265 52.795 201.435 ;
        RECT 53.585 201.265 53.755 201.435 ;
        RECT 54.045 201.265 54.215 201.435 ;
        RECT 54.505 201.265 54.675 201.435 ;
        RECT 54.965 201.265 55.135 201.435 ;
        RECT 55.425 201.265 55.595 201.435 ;
        RECT 55.885 201.265 56.055 201.435 ;
        RECT 56.345 201.265 56.515 201.435 ;
        RECT 57.335 201.265 57.505 201.435 ;
        RECT 58.335 201.265 58.505 201.435 ;
        RECT 58.795 201.265 58.965 201.435 ;
        RECT 59.255 201.265 59.425 201.435 ;
        RECT 59.715 201.265 59.885 201.435 ;
        RECT 60.175 201.265 60.345 201.435 ;
        RECT 61.135 201.265 61.305 201.435 ;
        RECT 61.595 201.265 61.765 201.435 ;
        RECT 62.055 201.265 62.225 201.435 ;
        RECT 62.515 201.265 62.685 201.435 ;
        RECT 62.975 201.265 63.145 201.435 ;
        RECT 63.435 201.265 63.605 201.435 ;
        RECT 63.895 201.265 64.065 201.435 ;
        RECT 64.885 201.265 65.055 201.435 ;
        RECT 65.345 201.265 65.515 201.435 ;
        RECT 65.805 201.265 65.975 201.435 ;
        RECT 66.265 201.265 66.435 201.435 ;
        RECT 66.725 201.265 66.895 201.435 ;
        RECT 67.685 201.265 67.855 201.435 ;
        RECT 68.145 201.265 68.315 201.435 ;
        RECT 68.605 201.265 68.775 201.435 ;
        RECT 69.065 201.265 69.235 201.435 ;
        RECT 69.525 201.265 69.695 201.435 ;
        RECT 69.985 201.265 70.155 201.435 ;
        RECT 70.445 201.265 70.615 201.435 ;
        RECT 71.445 201.265 71.615 201.435 ;
        RECT 72.495 201.265 72.665 201.435 ;
        RECT 72.955 201.265 73.125 201.435 ;
        RECT 73.415 201.265 73.585 201.435 ;
        RECT 73.875 201.265 74.045 201.435 ;
        RECT 74.335 201.265 74.505 201.435 ;
        RECT 75.395 201.265 75.565 201.435 ;
        RECT 75.855 201.265 76.025 201.435 ;
        RECT 76.315 201.265 76.485 201.435 ;
        RECT 76.775 201.265 76.945 201.435 ;
        RECT 77.235 201.265 77.405 201.435 ;
        RECT 77.695 201.265 77.865 201.435 ;
        RECT 78.155 201.265 78.325 201.435 ;
        RECT 30.945 200.625 31.115 200.795 ;
        RECT 31.405 200.625 31.575 200.795 ;
        RECT 31.865 200.625 32.035 200.795 ;
        RECT 32.325 200.625 32.495 200.795 ;
        RECT 32.785 200.625 32.955 200.795 ;
        RECT 33.245 200.625 33.415 200.795 ;
        RECT 34.045 200.625 34.215 200.795 ;
        RECT 34.505 200.625 34.675 200.795 ;
        RECT 34.965 200.625 35.135 200.795 ;
        RECT 35.425 200.625 35.595 200.795 ;
        RECT 35.885 200.625 36.055 200.795 ;
        RECT 36.345 200.625 36.515 200.795 ;
        RECT 37.015 200.635 37.185 200.805 ;
        RECT 37.475 200.635 37.645 200.805 ;
        RECT 37.935 200.635 38.105 200.805 ;
        RECT 38.395 200.635 38.565 200.805 ;
        RECT 38.855 200.635 39.025 200.805 ;
        RECT 39.315 200.635 39.485 200.805 ;
        RECT 40.145 200.635 40.315 200.805 ;
        RECT 40.605 200.635 40.775 200.805 ;
        RECT 41.065 200.635 41.235 200.805 ;
        RECT 41.525 200.635 41.695 200.805 ;
        RECT 41.985 200.635 42.155 200.805 ;
        RECT 42.445 200.635 42.615 200.805 ;
        RECT 43.185 200.635 43.355 200.805 ;
        RECT 44.235 200.635 44.405 200.805 ;
        RECT 44.695 200.635 44.865 200.805 ;
        RECT 45.155 200.635 45.325 200.805 ;
        RECT 45.615 200.635 45.785 200.805 ;
        RECT 46.075 200.635 46.245 200.805 ;
        RECT 46.535 200.635 46.705 200.805 ;
        RECT 47.395 200.635 47.565 200.805 ;
        RECT 47.855 200.635 48.025 200.805 ;
        RECT 48.315 200.635 48.485 200.805 ;
        RECT 48.775 200.635 48.945 200.805 ;
        RECT 49.235 200.635 49.405 200.805 ;
        RECT 49.695 200.635 49.865 200.805 ;
        RECT 50.785 200.635 50.955 200.805 ;
        RECT 51.245 200.635 51.415 200.805 ;
        RECT 51.705 200.635 51.875 200.805 ;
        RECT 52.165 200.635 52.335 200.805 ;
        RECT 52.625 200.635 52.795 200.805 ;
        RECT 53.085 200.635 53.255 200.805 ;
        RECT 53.945 200.635 54.115 200.805 ;
        RECT 54.405 200.635 54.575 200.805 ;
        RECT 54.865 200.635 55.035 200.805 ;
        RECT 55.325 200.635 55.495 200.805 ;
        RECT 55.785 200.635 55.955 200.805 ;
        RECT 56.245 200.635 56.415 200.805 ;
        RECT 57.335 200.645 57.505 200.815 ;
        RECT 58.335 200.645 58.505 200.815 ;
        RECT 58.795 200.645 58.965 200.815 ;
        RECT 59.255 200.645 59.425 200.815 ;
        RECT 59.715 200.645 59.885 200.815 ;
        RECT 60.175 200.645 60.345 200.815 ;
        RECT 60.635 200.645 60.805 200.815 ;
        RECT 61.535 200.645 61.705 200.815 ;
        RECT 61.995 200.645 62.165 200.815 ;
        RECT 62.455 200.645 62.625 200.815 ;
        RECT 62.915 200.645 63.085 200.815 ;
        RECT 63.375 200.645 63.545 200.815 ;
        RECT 63.835 200.645 64.005 200.815 ;
        RECT 64.885 200.645 65.055 200.815 ;
        RECT 65.345 200.645 65.515 200.815 ;
        RECT 65.805 200.645 65.975 200.815 ;
        RECT 66.265 200.645 66.435 200.815 ;
        RECT 66.725 200.645 66.895 200.815 ;
        RECT 67.185 200.645 67.355 200.815 ;
        RECT 68.085 200.645 68.255 200.815 ;
        RECT 68.545 200.645 68.715 200.815 ;
        RECT 69.005 200.645 69.175 200.815 ;
        RECT 69.465 200.645 69.635 200.815 ;
        RECT 69.925 200.645 70.095 200.815 ;
        RECT 70.385 200.645 70.555 200.815 ;
        RECT 71.445 200.645 71.615 200.815 ;
        RECT 72.495 200.645 72.665 200.815 ;
        RECT 72.955 200.645 73.125 200.815 ;
        RECT 73.415 200.645 73.585 200.815 ;
        RECT 73.875 200.645 74.045 200.815 ;
        RECT 74.335 200.645 74.505 200.815 ;
        RECT 74.795 200.645 74.965 200.815 ;
        RECT 75.855 200.645 76.025 200.815 ;
        RECT 76.315 200.645 76.485 200.815 ;
        RECT 76.775 200.645 76.945 200.815 ;
        RECT 77.235 200.645 77.405 200.815 ;
        RECT 77.695 200.645 77.865 200.815 ;
        RECT 78.155 200.645 78.325 200.815 ;
        RECT 30.985 200.070 31.155 200.250 ;
        RECT 31.865 199.065 32.090 199.265 ;
        RECT 33.200 199.065 33.370 199.235 ;
        RECT 37.055 198.475 37.225 198.645 ;
        RECT 37.990 199.075 38.160 199.245 ;
        RECT 38.625 199.075 38.800 199.245 ;
        RECT 39.270 199.075 39.440 199.245 ;
        RECT 44.200 198.550 44.400 198.750 ;
        RECT 45.210 199.085 45.380 199.255 ;
        RECT 46.490 199.075 46.660 199.245 ;
        RECT 50.770 200.050 50.970 200.250 ;
        RECT 46.075 198.450 46.250 198.635 ;
        RECT 51.760 199.075 51.930 199.245 ;
        RECT 53.040 199.075 53.210 199.245 ;
        RECT 58.300 199.400 58.500 199.600 ;
        RECT 52.600 198.500 52.800 198.700 ;
        RECT 59.250 199.100 59.450 199.310 ;
        RECT 59.900 199.050 60.100 199.250 ;
        RECT 60.590 199.085 60.760 199.255 ;
        RECT 64.850 198.500 65.050 198.700 ;
        RECT 65.900 199.100 66.100 199.300 ;
        RECT 66.500 199.100 66.700 199.300 ;
        RECT 67.140 199.085 67.310 199.255 ;
        RECT 72.470 199.900 72.650 200.095 ;
        RECT 73.500 199.100 73.700 199.300 ;
        RECT 74.750 199.085 74.920 199.255 ;
        RECT 74.330 198.515 74.505 198.685 ;
        RECT 30.945 197.905 31.115 198.075 ;
        RECT 31.405 197.905 31.575 198.075 ;
        RECT 31.865 197.905 32.035 198.075 ;
        RECT 32.325 197.905 32.495 198.075 ;
        RECT 32.785 197.905 32.955 198.075 ;
        RECT 33.245 197.905 33.415 198.075 ;
        RECT 34.045 197.905 34.215 198.075 ;
        RECT 34.505 197.905 34.675 198.075 ;
        RECT 34.965 197.905 35.135 198.075 ;
        RECT 35.425 197.905 35.595 198.075 ;
        RECT 35.885 197.905 36.055 198.075 ;
        RECT 36.345 197.905 36.515 198.075 ;
        RECT 37.015 197.915 37.185 198.085 ;
        RECT 37.475 197.915 37.645 198.085 ;
        RECT 37.935 197.915 38.105 198.085 ;
        RECT 38.395 197.915 38.565 198.085 ;
        RECT 38.855 197.915 39.025 198.085 ;
        RECT 39.315 197.915 39.485 198.085 ;
        RECT 40.145 197.915 40.315 198.085 ;
        RECT 40.605 197.915 40.775 198.085 ;
        RECT 41.065 197.915 41.235 198.085 ;
        RECT 41.525 197.915 41.695 198.085 ;
        RECT 41.985 197.915 42.155 198.085 ;
        RECT 42.445 197.915 42.615 198.085 ;
        RECT 43.185 197.915 43.355 198.085 ;
        RECT 44.235 197.915 44.405 198.085 ;
        RECT 44.695 197.915 44.865 198.085 ;
        RECT 45.155 197.915 45.325 198.085 ;
        RECT 45.615 197.915 45.785 198.085 ;
        RECT 46.075 197.915 46.245 198.085 ;
        RECT 46.535 197.915 46.705 198.085 ;
        RECT 47.395 197.915 47.565 198.085 ;
        RECT 47.855 197.915 48.025 198.085 ;
        RECT 48.315 197.915 48.485 198.085 ;
        RECT 48.775 197.915 48.945 198.085 ;
        RECT 49.235 197.915 49.405 198.085 ;
        RECT 49.695 197.915 49.865 198.085 ;
        RECT 50.785 197.915 50.955 198.085 ;
        RECT 51.245 197.915 51.415 198.085 ;
        RECT 51.705 197.915 51.875 198.085 ;
        RECT 52.165 197.915 52.335 198.085 ;
        RECT 52.625 197.915 52.795 198.085 ;
        RECT 53.085 197.915 53.255 198.085 ;
        RECT 53.945 197.915 54.115 198.085 ;
        RECT 54.405 197.915 54.575 198.085 ;
        RECT 54.865 197.915 55.035 198.085 ;
        RECT 55.325 197.915 55.495 198.085 ;
        RECT 55.785 197.915 55.955 198.085 ;
        RECT 56.245 197.915 56.415 198.085 ;
        RECT 57.335 197.925 57.505 198.095 ;
        RECT 58.335 197.925 58.505 198.095 ;
        RECT 58.795 197.925 58.965 198.095 ;
        RECT 59.255 197.925 59.425 198.095 ;
        RECT 59.715 197.925 59.885 198.095 ;
        RECT 60.175 197.925 60.345 198.095 ;
        RECT 60.635 197.925 60.805 198.095 ;
        RECT 61.535 197.925 61.705 198.095 ;
        RECT 61.995 197.925 62.165 198.095 ;
        RECT 62.455 197.925 62.625 198.095 ;
        RECT 62.915 197.925 63.085 198.095 ;
        RECT 63.375 197.925 63.545 198.095 ;
        RECT 63.835 197.925 64.005 198.095 ;
        RECT 64.885 197.925 65.055 198.095 ;
        RECT 65.345 197.925 65.515 198.095 ;
        RECT 65.805 197.925 65.975 198.095 ;
        RECT 66.265 197.925 66.435 198.095 ;
        RECT 66.725 197.925 66.895 198.095 ;
        RECT 67.185 197.925 67.355 198.095 ;
        RECT 68.085 197.925 68.255 198.095 ;
        RECT 68.545 197.925 68.715 198.095 ;
        RECT 69.005 197.925 69.175 198.095 ;
        RECT 69.465 197.925 69.635 198.095 ;
        RECT 69.925 197.925 70.095 198.095 ;
        RECT 70.385 197.925 70.555 198.095 ;
        RECT 71.445 197.925 71.615 198.095 ;
        RECT 72.495 197.925 72.665 198.095 ;
        RECT 72.955 197.925 73.125 198.095 ;
        RECT 73.415 197.925 73.585 198.095 ;
        RECT 73.875 197.925 74.045 198.095 ;
        RECT 74.335 197.925 74.505 198.095 ;
        RECT 74.795 197.925 74.965 198.095 ;
        RECT 75.855 197.925 76.025 198.095 ;
        RECT 76.315 197.925 76.485 198.095 ;
        RECT 76.775 197.925 76.945 198.095 ;
        RECT 77.235 197.925 77.405 198.095 ;
        RECT 77.695 197.925 77.865 198.095 ;
        RECT 78.155 197.925 78.325 198.095 ;
        RECT 30.945 197.275 31.115 197.445 ;
        RECT 31.405 197.275 31.575 197.445 ;
        RECT 31.865 197.275 32.035 197.445 ;
        RECT 32.325 197.275 32.495 197.445 ;
        RECT 32.785 197.275 32.955 197.445 ;
        RECT 33.245 197.275 33.415 197.445 ;
        RECT 33.705 197.275 33.875 197.445 ;
        RECT 34.585 197.275 34.755 197.445 ;
        RECT 35.045 197.275 35.215 197.445 ;
        RECT 35.505 197.275 35.675 197.445 ;
        RECT 35.965 197.275 36.135 197.445 ;
        RECT 37.015 197.275 37.185 197.445 ;
        RECT 37.475 197.275 37.645 197.445 ;
        RECT 37.935 197.275 38.105 197.445 ;
        RECT 38.395 197.275 38.565 197.445 ;
        RECT 38.855 197.275 39.025 197.445 ;
        RECT 39.315 197.275 39.485 197.445 ;
        RECT 39.775 197.275 39.945 197.445 ;
        RECT 40.805 197.275 40.975 197.445 ;
        RECT 41.265 197.275 41.435 197.445 ;
        RECT 41.725 197.275 41.895 197.445 ;
        RECT 42.185 197.275 42.355 197.445 ;
        RECT 43.185 197.275 43.355 197.445 ;
        RECT 44.235 197.275 44.405 197.445 ;
        RECT 44.695 197.275 44.865 197.445 ;
        RECT 45.155 197.275 45.325 197.445 ;
        RECT 45.615 197.275 45.785 197.445 ;
        RECT 46.075 197.275 46.245 197.445 ;
        RECT 46.535 197.275 46.705 197.445 ;
        RECT 46.995 197.275 47.165 197.445 ;
        RECT 47.745 197.275 47.915 197.445 ;
        RECT 48.205 197.275 48.375 197.445 ;
        RECT 48.665 197.275 48.835 197.445 ;
        RECT 49.125 197.275 49.295 197.445 ;
        RECT 49.585 197.275 49.755 197.445 ;
        RECT 50.045 197.275 50.215 197.445 ;
        RECT 50.785 197.275 50.955 197.445 ;
        RECT 51.245 197.275 51.415 197.445 ;
        RECT 51.705 197.275 51.875 197.445 ;
        RECT 52.165 197.275 52.335 197.445 ;
        RECT 52.625 197.275 52.795 197.445 ;
        RECT 53.085 197.275 53.255 197.445 ;
        RECT 53.545 197.275 53.715 197.445 ;
        RECT 54.385 197.275 54.555 197.445 ;
        RECT 54.845 197.275 55.015 197.445 ;
        RECT 55.305 197.275 55.475 197.445 ;
        RECT 55.765 197.275 55.935 197.445 ;
        RECT 56.225 197.275 56.395 197.445 ;
        RECT 56.685 197.275 56.855 197.445 ;
        RECT 57.335 197.275 57.505 197.445 ;
        RECT 58.335 197.275 58.505 197.445 ;
        RECT 58.795 197.275 58.965 197.445 ;
        RECT 59.255 197.275 59.425 197.445 ;
        RECT 59.715 197.275 59.885 197.445 ;
        RECT 60.175 197.275 60.345 197.445 ;
        RECT 60.635 197.275 60.805 197.445 ;
        RECT 61.095 197.275 61.265 197.445 ;
        RECT 62.035 197.275 62.205 197.445 ;
        RECT 62.495 197.275 62.665 197.445 ;
        RECT 62.955 197.275 63.125 197.445 ;
        RECT 63.415 197.275 63.585 197.445 ;
        RECT 63.875 197.275 64.045 197.445 ;
        RECT 64.335 197.275 64.505 197.445 ;
        RECT 64.885 197.275 65.055 197.445 ;
        RECT 65.345 197.275 65.515 197.445 ;
        RECT 65.805 197.275 65.975 197.445 ;
        RECT 66.265 197.275 66.435 197.445 ;
        RECT 66.725 197.275 66.895 197.445 ;
        RECT 67.185 197.275 67.355 197.445 ;
        RECT 67.645 197.275 67.815 197.445 ;
        RECT 68.535 197.275 68.705 197.445 ;
        RECT 68.995 197.275 69.165 197.445 ;
        RECT 69.455 197.275 69.625 197.445 ;
        RECT 69.915 197.275 70.085 197.445 ;
        RECT 70.375 197.275 70.545 197.445 ;
        RECT 70.835 197.275 71.005 197.445 ;
        RECT 71.445 197.275 71.615 197.445 ;
        RECT 72.485 197.275 72.655 197.445 ;
        RECT 72.945 197.275 73.115 197.445 ;
        RECT 73.405 197.275 73.575 197.445 ;
        RECT 73.865 197.275 74.035 197.445 ;
        RECT 74.325 197.275 74.495 197.445 ;
        RECT 74.785 197.275 74.955 197.445 ;
        RECT 75.245 197.275 75.415 197.445 ;
        RECT 76.775 197.275 76.945 197.445 ;
        RECT 77.235 197.275 77.405 197.445 ;
        RECT 77.695 197.275 77.865 197.445 ;
        RECT 78.155 197.275 78.325 197.445 ;
        RECT 33.650 196.500 33.850 196.700 ;
        RECT 31.225 195.715 31.395 195.885 ;
        RECT 31.810 195.715 32.010 195.915 ;
        RECT 39.705 196.515 39.875 196.685 ;
        RECT 37.300 195.650 37.500 195.900 ;
        RECT 37.880 195.715 38.050 195.885 ;
        RECT 44.535 195.700 44.715 195.885 ;
        RECT 45.100 195.715 45.270 195.885 ;
        RECT 46.995 196.085 47.165 196.255 ;
        RECT 51.065 195.715 51.235 195.885 ;
        RECT 51.650 195.715 51.820 195.885 ;
        RECT 53.500 196.050 53.700 196.250 ;
        RECT 58.615 195.715 58.785 195.885 ;
        RECT 59.200 195.715 59.370 195.885 ;
        RECT 61.050 196.100 61.250 196.300 ;
        RECT 65.165 195.715 65.335 195.885 ;
        RECT 65.750 195.715 65.920 195.885 ;
        RECT 67.245 195.200 67.415 195.385 ;
        RECT 72.800 196.000 72.975 196.170 ;
        RECT 73.350 195.715 73.520 195.885 ;
        RECT 75.250 196.100 75.450 196.300 ;
        RECT 30.945 194.555 31.115 194.725 ;
        RECT 31.405 194.555 31.575 194.725 ;
        RECT 31.865 194.555 32.035 194.725 ;
        RECT 32.325 194.555 32.495 194.725 ;
        RECT 32.785 194.555 32.955 194.725 ;
        RECT 33.245 194.555 33.415 194.725 ;
        RECT 33.705 194.555 33.875 194.725 ;
        RECT 34.585 194.555 34.755 194.725 ;
        RECT 35.045 194.555 35.215 194.725 ;
        RECT 35.505 194.555 35.675 194.725 ;
        RECT 35.965 194.555 36.135 194.725 ;
        RECT 37.015 194.555 37.185 194.725 ;
        RECT 37.475 194.555 37.645 194.725 ;
        RECT 37.935 194.555 38.105 194.725 ;
        RECT 38.395 194.555 38.565 194.725 ;
        RECT 38.855 194.555 39.025 194.725 ;
        RECT 39.315 194.555 39.485 194.725 ;
        RECT 39.775 194.555 39.945 194.725 ;
        RECT 40.805 194.555 40.975 194.725 ;
        RECT 41.265 194.555 41.435 194.725 ;
        RECT 41.725 194.555 41.895 194.725 ;
        RECT 42.185 194.555 42.355 194.725 ;
        RECT 43.185 194.555 43.355 194.725 ;
        RECT 44.235 194.555 44.405 194.725 ;
        RECT 44.695 194.555 44.865 194.725 ;
        RECT 45.155 194.555 45.325 194.725 ;
        RECT 45.615 194.555 45.785 194.725 ;
        RECT 46.075 194.555 46.245 194.725 ;
        RECT 46.535 194.555 46.705 194.725 ;
        RECT 46.995 194.555 47.165 194.725 ;
        RECT 47.745 194.555 47.915 194.725 ;
        RECT 48.205 194.555 48.375 194.725 ;
        RECT 48.665 194.555 48.835 194.725 ;
        RECT 49.125 194.555 49.295 194.725 ;
        RECT 49.585 194.555 49.755 194.725 ;
        RECT 50.045 194.555 50.215 194.725 ;
        RECT 50.785 194.555 50.955 194.725 ;
        RECT 51.245 194.555 51.415 194.725 ;
        RECT 51.705 194.555 51.875 194.725 ;
        RECT 52.165 194.555 52.335 194.725 ;
        RECT 52.625 194.555 52.795 194.725 ;
        RECT 53.085 194.555 53.255 194.725 ;
        RECT 53.545 194.555 53.715 194.725 ;
        RECT 54.385 194.555 54.555 194.725 ;
        RECT 54.845 194.555 55.015 194.725 ;
        RECT 55.305 194.555 55.475 194.725 ;
        RECT 55.765 194.555 55.935 194.725 ;
        RECT 56.225 194.555 56.395 194.725 ;
        RECT 56.685 194.555 56.855 194.725 ;
        RECT 57.335 194.555 57.505 194.725 ;
        RECT 58.335 194.555 58.505 194.725 ;
        RECT 58.795 194.555 58.965 194.725 ;
        RECT 59.255 194.555 59.425 194.725 ;
        RECT 59.715 194.555 59.885 194.725 ;
        RECT 60.175 194.555 60.345 194.725 ;
        RECT 60.635 194.555 60.805 194.725 ;
        RECT 61.095 194.555 61.265 194.725 ;
        RECT 62.035 194.555 62.205 194.725 ;
        RECT 62.495 194.555 62.665 194.725 ;
        RECT 62.955 194.555 63.125 194.725 ;
        RECT 63.415 194.555 63.585 194.725 ;
        RECT 63.875 194.555 64.045 194.725 ;
        RECT 64.335 194.555 64.505 194.725 ;
        RECT 64.885 194.555 65.055 194.725 ;
        RECT 65.345 194.555 65.515 194.725 ;
        RECT 65.805 194.555 65.975 194.725 ;
        RECT 66.265 194.555 66.435 194.725 ;
        RECT 66.725 194.555 66.895 194.725 ;
        RECT 67.185 194.555 67.355 194.725 ;
        RECT 67.645 194.555 67.815 194.725 ;
        RECT 68.535 194.555 68.705 194.725 ;
        RECT 68.995 194.555 69.165 194.725 ;
        RECT 69.455 194.555 69.625 194.725 ;
        RECT 69.915 194.555 70.085 194.725 ;
        RECT 70.375 194.555 70.545 194.725 ;
        RECT 70.835 194.555 71.005 194.725 ;
        RECT 71.445 194.555 71.615 194.725 ;
        RECT 72.485 194.555 72.655 194.725 ;
        RECT 72.945 194.555 73.115 194.725 ;
        RECT 73.405 194.555 73.575 194.725 ;
        RECT 73.865 194.555 74.035 194.725 ;
        RECT 74.325 194.555 74.495 194.725 ;
        RECT 74.785 194.555 74.955 194.725 ;
        RECT 75.245 194.555 75.415 194.725 ;
        RECT 76.775 194.555 76.945 194.725 ;
        RECT 77.235 194.555 77.405 194.725 ;
        RECT 77.695 194.555 77.865 194.725 ;
        RECT 78.155 194.555 78.325 194.725 ;
      LAYER met1 ;
        RECT 30.800 203.830 78.470 204.310 ;
        RECT 74.050 203.200 74.500 203.650 ;
        RECT 30.850 202.450 31.250 202.850 ;
        RECT 31.750 202.400 32.150 202.800 ;
        RECT 33.450 202.650 33.895 203.000 ;
        RECT 34.100 202.700 34.500 202.800 ;
        RECT 33.450 202.600 33.850 202.650 ;
        RECT 34.050 202.400 34.600 202.700 ;
        RECT 36.000 202.650 36.400 203.050 ;
        RECT 36.800 202.400 37.350 202.800 ;
        RECT 32.600 201.950 33.055 202.350 ;
        RECT 37.865 202.300 38.250 202.700 ;
        RECT 40.300 202.350 40.700 202.750 ;
        RECT 42.150 202.700 42.550 203.100 ;
        RECT 40.930 202.600 41.300 202.640 ;
        RECT 38.750 201.950 39.150 202.350 ;
        RECT 40.900 202.200 41.300 202.600 ;
        RECT 44.200 202.350 44.600 202.750 ;
        RECT 45.050 202.300 45.450 202.750 ;
        RECT 46.050 202.300 46.450 202.700 ;
        RECT 47.365 202.650 47.610 202.700 ;
        RECT 47.200 202.345 47.610 202.650 ;
        RECT 47.850 202.350 48.250 202.750 ;
        RECT 49.700 202.700 50.100 203.100 ;
        RECT 56.150 202.750 56.550 203.150 ;
        RECT 50.600 202.350 51.000 202.750 ;
        RECT 51.635 202.650 51.975 202.675 ;
        RECT 47.200 202.300 47.600 202.345 ;
        RECT 51.600 202.250 52.000 202.650 ;
        RECT 52.600 202.250 53.000 202.650 ;
        RECT 54.300 202.350 54.800 202.700 ;
        RECT 55.000 202.245 55.400 202.705 ;
        RECT 58.250 202.400 58.650 202.800 ;
        RECT 59.150 202.200 59.600 202.750 ;
        RECT 60.100 202.550 60.500 202.950 ;
        RECT 63.700 202.750 64.100 203.150 ;
        RECT 61.800 202.200 62.450 202.650 ;
        RECT 62.600 202.250 63.000 202.650 ;
        RECT 64.700 202.300 65.100 202.700 ;
        RECT 65.700 202.300 66.100 202.700 ;
        RECT 68.400 202.650 68.800 202.750 ;
        RECT 70.300 202.650 70.700 203.050 ;
        RECT 72.250 202.700 72.700 202.900 ;
        RECT 66.650 202.250 67.050 202.650 ;
        RECT 67.795 202.200 68.200 202.650 ;
        RECT 68.350 202.400 68.950 202.650 ;
        RECT 72.250 202.400 72.795 202.700 ;
        RECT 68.400 202.350 68.800 202.400 ;
        RECT 73.300 202.300 73.750 202.700 ;
        RECT 76.050 202.300 76.700 202.700 ;
        RECT 76.850 202.300 77.350 202.750 ;
        RECT 78.000 202.700 78.400 203.100 ;
        RECT 30.800 201.110 78.470 201.590 ;
        RECT 33.035 201.105 33.390 201.110 ;
        RECT 36.370 201.105 36.915 201.110 ;
        RECT 42.560 201.105 43.105 201.110 ;
        RECT 57.190 200.960 78.470 200.970 ;
        RECT 36.870 200.950 78.470 200.960 ;
        RECT 30.800 200.490 78.470 200.950 ;
        RECT 30.800 200.480 56.560 200.490 ;
        RECT 30.800 200.470 36.660 200.480 ;
        RECT 30.900 199.900 31.300 200.300 ;
        RECT 50.700 199.900 51.100 200.300 ;
        RECT 72.350 199.850 72.750 200.250 ;
        RECT 31.700 199.350 32.100 199.400 ;
        RECT 31.700 199.000 32.150 199.350 ;
        RECT 33.150 199.000 33.550 199.400 ;
        RECT 37.900 199.325 38.300 199.400 ;
        RECT 37.885 199.010 38.345 199.325 ;
        RECT 37.900 199.000 38.300 199.010 ;
        RECT 38.550 199.000 38.950 199.450 ;
        RECT 39.200 199.000 39.600 199.400 ;
        RECT 45.050 199.050 45.450 199.450 ;
        RECT 46.450 199.000 46.850 199.400 ;
        RECT 51.650 199.000 52.050 199.400 ;
        RECT 53.000 199.000 53.400 199.400 ;
        RECT 58.200 199.300 58.600 199.700 ;
        RECT 59.150 199.050 59.550 199.450 ;
        RECT 59.800 199.000 60.200 199.400 ;
        RECT 60.500 199.000 60.900 199.400 ;
        RECT 65.750 199.000 66.150 199.400 ;
        RECT 66.400 199.000 66.800 199.400 ;
        RECT 67.100 199.000 67.500 199.400 ;
        RECT 73.400 199.000 73.800 199.400 ;
        RECT 74.700 198.950 75.100 199.350 ;
        RECT 32.700 198.400 33.100 198.800 ;
        RECT 36.900 198.400 37.300 198.800 ;
        RECT 44.050 198.450 44.450 198.850 ;
        RECT 45.950 198.400 46.350 198.800 ;
        RECT 52.450 198.400 52.850 198.800 ;
        RECT 64.700 198.400 65.100 198.800 ;
        RECT 74.150 198.450 74.550 198.850 ;
        RECT 56.520 198.240 78.470 198.250 ;
        RECT 36.870 198.230 78.470 198.240 ;
        RECT 30.800 197.770 78.470 198.230 ;
        RECT 30.800 197.760 57.215 197.770 ;
        RECT 30.800 197.750 36.660 197.760 ;
        RECT 56.520 197.750 57.215 197.760 ;
        RECT 30.800 197.120 78.470 197.600 ;
        RECT 33.600 196.400 34.000 196.800 ;
        RECT 39.650 196.400 40.050 196.800 ;
        RECT 31.095 195.600 31.500 196.000 ;
        RECT 31.700 195.650 32.100 196.050 ;
        RECT 37.200 195.550 37.600 195.950 ;
        RECT 37.800 195.600 38.200 196.000 ;
        RECT 44.400 195.600 44.800 196.000 ;
        RECT 45.000 195.650 45.400 196.050 ;
        RECT 46.900 196.000 47.300 196.400 ;
        RECT 50.900 195.650 51.300 196.050 ;
        RECT 51.550 195.650 51.950 196.050 ;
        RECT 53.400 196.000 53.800 196.400 ;
        RECT 58.500 195.600 58.900 196.000 ;
        RECT 59.150 195.650 59.550 196.050 ;
        RECT 60.950 196.000 61.400 196.800 ;
        RECT 65.050 195.600 65.450 196.000 ;
        RECT 65.650 195.600 66.050 196.000 ;
        RECT 72.650 195.950 73.050 196.350 ;
        RECT 73.250 195.650 73.650 196.050 ;
        RECT 75.150 196.000 75.550 196.400 ;
        RECT 67.150 195.150 67.600 195.550 ;
        RECT 67.150 195.100 67.345 195.150 ;
        RECT 30.800 194.400 78.470 194.880 ;
      LAYER via ;
        RECT 30.850 203.900 31.150 204.200 ;
        RECT 71.350 203.900 71.700 204.250 ;
        RECT 74.100 203.250 74.450 203.600 ;
        RECT 30.900 202.500 31.200 202.800 ;
        RECT 31.800 202.400 32.100 202.710 ;
        RECT 33.500 202.650 33.800 202.950 ;
        RECT 34.150 202.450 34.450 202.750 ;
        RECT 36.050 202.700 36.350 203.000 ;
        RECT 42.200 202.750 42.500 203.050 ;
        RECT 49.750 202.750 50.050 203.050 ;
        RECT 56.200 202.800 56.500 203.100 ;
        RECT 36.850 202.450 37.150 202.750 ;
        RECT 37.900 202.350 38.200 202.650 ;
        RECT 40.350 202.400 40.650 202.700 ;
        RECT 32.700 202.000 33.000 202.300 ;
        RECT 38.800 202.000 39.100 202.300 ;
        RECT 40.950 202.250 41.250 202.550 ;
        RECT 44.250 202.400 44.550 202.700 ;
        RECT 45.100 202.400 45.400 202.700 ;
        RECT 46.100 202.350 46.400 202.650 ;
        RECT 47.250 202.300 47.550 202.600 ;
        RECT 47.900 202.400 48.200 202.700 ;
        RECT 50.650 202.400 50.950 202.700 ;
        RECT 51.650 202.300 51.950 202.600 ;
        RECT 52.650 202.300 52.950 202.600 ;
        RECT 54.400 202.400 54.700 202.700 ;
        RECT 55.050 202.345 55.350 202.650 ;
        RECT 58.300 202.450 58.600 202.750 ;
        RECT 59.200 202.400 59.500 202.700 ;
        RECT 60.150 202.600 60.450 202.900 ;
        RECT 63.750 202.800 64.050 203.100 ;
        RECT 61.900 202.300 62.200 202.600 ;
        RECT 62.650 202.300 62.950 202.600 ;
        RECT 64.750 202.350 65.050 202.650 ;
        RECT 65.750 202.350 66.050 202.650 ;
        RECT 66.700 202.300 67.000 202.600 ;
        RECT 67.850 202.300 68.150 202.600 ;
        RECT 68.450 202.400 68.750 202.700 ;
        RECT 70.350 202.700 70.650 203.000 ;
        RECT 72.300 202.500 72.600 202.800 ;
        RECT 78.050 202.750 78.350 203.050 ;
        RECT 73.350 202.350 73.650 202.650 ;
        RECT 76.100 202.350 76.400 202.650 ;
        RECT 76.900 202.350 77.200 202.650 ;
        RECT 57.250 201.200 57.600 201.550 ;
        RECT 71.350 200.500 71.700 200.850 ;
        RECT 30.950 199.950 31.250 200.250 ;
        RECT 50.750 199.950 51.050 200.250 ;
        RECT 72.400 199.900 72.700 200.200 ;
        RECT 31.750 199.050 32.050 199.350 ;
        RECT 33.200 199.050 33.500 199.350 ;
        RECT 37.950 199.050 38.250 199.350 ;
        RECT 38.600 199.050 38.900 199.350 ;
        RECT 39.250 199.050 39.550 199.350 ;
        RECT 45.100 199.100 45.400 199.400 ;
        RECT 46.500 199.050 46.800 199.350 ;
        RECT 51.700 199.050 52.000 199.350 ;
        RECT 53.050 199.050 53.350 199.350 ;
        RECT 58.250 199.350 58.550 199.650 ;
        RECT 59.200 199.100 59.500 199.400 ;
        RECT 59.850 199.050 60.150 199.350 ;
        RECT 60.550 199.050 60.850 199.355 ;
        RECT 65.800 199.050 66.100 199.350 ;
        RECT 66.450 199.050 66.750 199.350 ;
        RECT 67.150 199.050 67.450 199.350 ;
        RECT 73.450 199.050 73.750 199.350 ;
        RECT 74.750 199.000 75.050 199.300 ;
        RECT 32.750 198.450 33.050 198.750 ;
        RECT 36.950 198.450 37.250 198.750 ;
        RECT 44.100 198.500 44.400 198.800 ;
        RECT 46.000 198.450 46.300 198.750 ;
        RECT 52.500 198.450 52.800 198.750 ;
        RECT 64.750 198.450 65.050 198.750 ;
        RECT 74.200 198.500 74.500 198.800 ;
        RECT 57.250 197.850 57.600 198.200 ;
        RECT 71.350 197.150 71.700 197.500 ;
        RECT 33.650 196.450 33.950 196.750 ;
        RECT 39.695 196.450 39.995 196.750 ;
        RECT 61.050 196.500 61.350 196.800 ;
        RECT 46.950 196.050 47.250 196.350 ;
        RECT 53.450 196.050 53.750 196.350 ;
        RECT 31.150 195.650 31.450 195.950 ;
        RECT 31.750 195.700 32.050 196.000 ;
        RECT 37.250 195.600 37.550 195.910 ;
        RECT 37.850 195.650 38.150 195.950 ;
        RECT 44.450 195.650 44.750 195.950 ;
        RECT 45.050 195.700 45.350 196.000 ;
        RECT 50.950 195.700 51.250 196.000 ;
        RECT 72.700 196.000 73.000 196.300 ;
        RECT 75.200 196.050 75.500 196.350 ;
        RECT 51.600 195.700 51.900 196.000 ;
        RECT 58.550 195.650 58.850 195.950 ;
        RECT 59.200 195.700 59.500 196.000 ;
        RECT 65.100 195.650 65.400 195.950 ;
        RECT 65.700 195.650 66.000 195.950 ;
        RECT 73.300 195.700 73.600 196.000 ;
        RECT 67.250 195.200 67.550 195.500 ;
        RECT 30.850 194.500 31.150 194.800 ;
        RECT 57.250 194.500 57.600 194.850 ;
      LAYER met2 ;
        RECT 30.100 203.800 31.200 204.300 ;
        RECT 30.800 203.150 31.300 203.650 ;
        RECT 30.850 202.450 31.250 203.150 ;
        RECT 31.750 202.250 32.150 202.800 ;
        RECT 33.450 202.600 33.950 203.000 ;
        RECT 31.700 201.750 32.150 202.250 ;
        RECT 32.600 201.950 33.050 202.350 ;
        RECT 33.550 202.250 33.950 202.600 ;
        RECT 34.100 202.400 34.500 203.650 ;
        RECT 36.750 203.150 37.200 203.650 ;
        RECT 36.000 202.650 36.400 203.050 ;
        RECT 36.800 202.400 37.200 203.150 ;
        RECT 40.300 202.800 40.750 203.650 ;
        RECT 32.700 201.450 33.000 201.950 ;
        RECT 33.500 201.750 33.950 202.250 ;
        RECT 37.865 202.200 38.250 202.700 ;
        RECT 37.750 201.700 38.250 202.200 ;
        RECT 31.700 201.050 32.100 201.450 ;
        RECT 32.600 201.050 33.000 201.450 ;
        RECT 30.900 199.900 31.300 200.300 ;
        RECT 31.700 199.500 32.000 201.050 ;
        RECT 31.700 199.010 32.100 199.500 ;
        RECT 33.150 199.350 33.550 199.400 ;
        RECT 33.100 199.000 33.550 199.350 ;
        RECT 37.900 199.000 38.300 201.100 ;
        RECT 38.750 200.700 39.150 202.350 ;
        RECT 40.250 202.300 40.750 202.800 ;
        RECT 42.150 202.700 42.550 203.100 ;
        RECT 40.900 201.695 41.300 202.600 ;
        RECT 44.200 202.350 44.600 204.000 ;
        RECT 45.050 201.450 45.450 202.745 ;
        RECT 46.000 202.250 46.500 202.750 ;
        RECT 47.200 201.450 47.600 202.650 ;
        RECT 47.850 202.350 48.250 204.000 ;
        RECT 49.700 202.700 50.100 203.100 ;
        RECT 50.600 202.350 51.000 203.600 ;
        RECT 54.400 202.700 54.800 203.500 ;
        RECT 56.150 202.750 56.550 203.150 ;
        RECT 51.600 202.405 52.000 202.650 ;
        RECT 51.600 201.545 52.005 202.405 ;
        RECT 38.550 199.950 38.950 200.350 ;
        RECT 44.900 200.150 45.400 200.250 ;
        RECT 38.600 199.450 38.900 199.950 ;
        RECT 44.900 199.750 45.450 200.150 ;
        RECT 50.700 199.900 51.100 200.300 ;
        RECT 38.550 199.000 38.950 199.450 ;
        RECT 39.200 199.000 39.600 199.400 ;
        RECT 45.050 199.050 45.450 199.750 ;
        RECT 33.100 198.950 33.500 199.000 ;
        RECT 46.400 198.950 46.900 199.450 ;
        RECT 51.650 199.000 52.050 201.250 ;
        RECT 52.600 200.850 53.000 202.650 ;
        RECT 54.300 202.350 54.800 202.700 ;
        RECT 54.995 202.050 55.400 202.695 ;
        RECT 58.250 202.400 58.650 203.750 ;
        RECT 61.550 203.200 62.300 203.750 ;
        RECT 54.850 201.550 55.400 202.050 ;
        RECT 59.150 202.000 59.550 202.750 ;
        RECT 60.100 202.550 60.500 202.950 ;
        RECT 61.900 202.650 62.300 203.200 ;
        RECT 63.700 202.750 64.100 203.150 ;
        RECT 61.750 202.200 62.450 202.650 ;
        RECT 62.600 202.000 63.000 202.650 ;
        RECT 64.700 202.300 65.100 203.700 ;
        RECT 54.850 201.545 55.000 201.550 ;
        RECT 53.000 199.000 53.400 199.400 ;
        RECT 32.700 198.150 33.150 198.800 ;
        RECT 36.900 198.200 37.300 198.800 ;
        RECT 44.050 197.450 44.450 198.860 ;
        RECT 45.950 198.250 46.350 198.800 ;
        RECT 34.900 196.800 35.300 197.000 ;
        RECT 40.900 196.800 41.400 196.900 ;
        RECT 31.100 195.600 31.500 196.650 ;
        RECT 33.600 196.400 35.300 196.800 ;
        RECT 39.645 196.400 41.400 196.800 ;
        RECT 44.400 196.400 44.900 196.900 ;
        RECT 31.700 195.400 32.100 196.050 ;
        RECT 37.200 195.550 37.600 195.950 ;
        RECT 37.750 195.550 38.250 196.050 ;
        RECT 44.400 195.600 44.800 196.400 ;
        RECT 44.950 195.600 45.450 196.100 ;
        RECT 46.900 196.000 49.250 196.400 ;
        RECT 52.450 196.050 52.850 198.800 ;
        RECT 48.850 195.650 49.250 196.000 ;
        RECT 37.250 195.250 37.550 195.550 ;
        RECT 50.900 195.300 51.300 196.050 ;
        RECT 51.550 195.650 52.850 196.050 ;
        RECT 53.400 196.000 55.000 196.400 ;
        RECT 37.250 195.150 37.650 195.250 ;
        RECT 30.800 194.400 31.200 194.900 ;
        RECT 37.250 194.650 37.750 195.150 ;
        RECT 50.850 194.800 51.350 195.300 ;
        RECT 57.200 194.400 57.650 201.600 ;
        RECT 59.150 201.500 59.750 202.000 ;
        RECT 62.495 201.500 63.000 202.000 ;
        RECT 65.700 201.450 66.095 202.700 ;
        RECT 66.650 202.250 67.050 202.650 ;
        RECT 67.795 202.200 68.200 202.650 ;
        RECT 68.400 202.350 68.800 203.700 ;
        RECT 70.300 202.650 70.700 203.050 ;
        RECT 67.800 201.950 68.200 202.200 ;
        RECT 67.700 201.450 68.250 201.950 ;
        RECT 58.200 200.500 58.600 201.000 ;
        RECT 66.350 200.500 66.800 201.000 ;
        RECT 58.200 199.700 58.550 200.500 ;
        RECT 58.200 199.300 58.600 199.700 ;
        RECT 58.500 195.600 58.900 198.100 ;
        RECT 59.150 196.650 59.550 199.450 ;
        RECT 59.800 197.700 60.200 200.300 ;
        RECT 60.500 199.000 60.900 199.400 ;
        RECT 65.750 199.000 66.150 200.150 ;
        RECT 66.400 199.000 66.800 200.500 ;
        RECT 67.100 199.000 67.500 199.400 ;
        RECT 64.700 198.300 65.100 198.800 ;
        RECT 71.300 197.050 71.750 204.300 ;
        RECT 72.250 202.400 72.700 203.900 ;
        RECT 74.050 203.200 74.500 203.650 ;
        RECT 75.950 203.400 76.450 203.900 ;
        RECT 73.300 202.250 73.700 202.700 ;
        RECT 73.200 201.600 73.700 202.250 ;
        RECT 72.350 199.850 72.750 201.200 ;
        RECT 73.400 199.000 73.800 200.450 ;
        RECT 74.050 200.050 74.450 203.200 ;
        RECT 76.050 202.300 76.450 203.400 ;
        RECT 76.850 202.300 77.350 202.750 ;
        RECT 78.000 202.700 78.400 203.100 ;
        RECT 76.850 202.150 77.250 202.300 ;
        RECT 76.750 201.600 77.250 202.150 ;
        RECT 74.700 198.950 75.100 199.750 ;
        RECT 62.600 196.850 63.100 196.950 ;
        RECT 60.950 196.450 63.100 196.850 ;
        RECT 59.150 195.650 59.550 196.050 ;
        RECT 65.050 195.600 65.450 196.850 ;
        RECT 65.650 195.600 66.050 196.000 ;
        RECT 72.650 195.950 73.050 198.650 ;
        RECT 74.150 198.450 74.550 198.850 ;
        RECT 67.200 195.150 69.800 195.550 ;
        RECT 73.250 194.950 73.650 196.050 ;
        RECT 75.150 196.000 76.400 196.400 ;
      LAYER via2 ;
        RECT 30.150 203.900 30.450 204.200 ;
        RECT 30.900 203.250 31.200 203.550 ;
        RECT 34.100 203.250 34.400 203.550 ;
        RECT 31.750 201.850 32.050 202.150 ;
        RECT 36.850 203.250 37.150 203.550 ;
        RECT 36.050 202.700 36.350 203.000 ;
        RECT 40.350 203.200 40.650 203.500 ;
        RECT 44.250 203.550 44.550 203.850 ;
        RECT 33.600 201.850 33.900 202.150 ;
        RECT 37.850 201.800 38.150 202.100 ;
        RECT 31.750 201.100 32.050 201.400 ;
        RECT 32.650 201.100 32.950 201.400 ;
        RECT 30.950 199.950 31.250 200.250 ;
        RECT 37.950 200.750 38.250 201.050 ;
        RECT 33.150 199.050 33.450 199.350 ;
        RECT 42.200 202.750 42.500 203.050 ;
        RECT 47.900 203.550 48.200 203.850 ;
        RECT 40.900 201.750 41.200 202.055 ;
        RECT 46.050 202.300 46.450 202.700 ;
        RECT 45.100 201.550 45.400 201.850 ;
        RECT 50.650 203.200 50.950 203.500 ;
        RECT 49.750 202.750 50.050 203.050 ;
        RECT 54.450 203.150 54.750 203.450 ;
        RECT 58.350 203.350 58.650 203.650 ;
        RECT 56.200 202.800 56.500 203.095 ;
        RECT 47.250 201.550 47.550 201.850 ;
        RECT 51.650 201.650 51.950 201.955 ;
        RECT 38.800 200.750 39.100 201.050 ;
        RECT 51.700 200.900 52.000 201.200 ;
        RECT 38.600 200.000 38.900 200.300 ;
        RECT 44.950 199.800 45.350 200.200 ;
        RECT 50.750 199.950 51.050 200.250 ;
        RECT 39.250 199.050 39.550 199.350 ;
        RECT 46.450 199.000 46.850 199.400 ;
        RECT 61.900 203.300 62.200 203.600 ;
        RECT 55.000 201.650 55.300 201.945 ;
        RECT 60.150 202.600 60.450 202.900 ;
        RECT 64.750 203.300 65.050 203.600 ;
        RECT 63.750 202.800 64.050 203.100 ;
        RECT 68.450 203.250 68.750 203.550 ;
        RECT 59.250 201.650 59.550 201.950 ;
        RECT 52.650 200.900 52.950 201.200 ;
        RECT 53.050 199.050 53.350 199.350 ;
        RECT 32.800 198.200 33.100 198.500 ;
        RECT 36.950 198.250 37.250 198.550 ;
        RECT 46.000 198.250 46.300 198.550 ;
        RECT 44.100 197.500 44.400 197.800 ;
        RECT 52.500 197.500 52.800 197.800 ;
        RECT 31.150 196.300 31.450 196.600 ;
        RECT 34.950 196.450 35.250 196.750 ;
        RECT 41.000 196.500 41.300 196.800 ;
        RECT 44.450 196.450 44.850 196.850 ;
        RECT 31.750 195.450 32.050 195.750 ;
        RECT 37.800 195.600 38.200 196.000 ;
        RECT 45.000 195.650 45.400 196.050 ;
        RECT 48.900 195.700 49.200 196.000 ;
        RECT 54.650 196.050 54.950 196.350 ;
        RECT 30.850 194.500 31.150 194.800 ;
        RECT 37.300 194.700 37.700 195.100 ;
        RECT 50.900 194.850 51.300 195.250 ;
        RECT 62.650 201.550 62.950 201.850 ;
        RECT 66.700 202.300 67.000 202.600 ;
        RECT 70.350 202.700 70.650 203.000 ;
        RECT 65.750 201.500 66.050 201.800 ;
        RECT 67.850 201.550 68.150 201.850 ;
        RECT 58.250 200.650 58.550 200.950 ;
        RECT 66.400 200.650 66.700 200.950 ;
        RECT 59.850 199.950 60.150 200.250 ;
        RECT 58.550 197.750 58.850 198.050 ;
        RECT 65.800 199.800 66.100 200.100 ;
        RECT 60.550 199.050 60.850 199.350 ;
        RECT 67.150 199.050 67.450 199.350 ;
        RECT 64.750 198.300 65.050 198.600 ;
        RECT 59.850 197.750 60.150 198.050 ;
        RECT 72.300 203.550 72.600 203.850 ;
        RECT 76.000 203.450 76.400 203.850 ;
        RECT 73.300 201.700 73.600 202.000 ;
        RECT 72.400 200.850 72.700 201.150 ;
        RECT 73.450 200.100 73.750 200.400 ;
        RECT 78.050 202.750 78.350 203.050 ;
        RECT 76.850 201.700 77.150 202.000 ;
        RECT 74.100 200.100 74.400 200.400 ;
        RECT 74.750 199.400 75.050 199.700 ;
        RECT 72.700 198.300 73.000 198.600 ;
        RECT 74.200 198.500 74.500 198.800 ;
        RECT 59.200 196.700 59.500 197.000 ;
        RECT 62.750 196.500 63.050 196.800 ;
        RECT 65.100 196.500 65.400 196.800 ;
        RECT 59.200 195.700 59.500 196.000 ;
        RECT 76.050 196.050 76.350 196.350 ;
        RECT 65.700 195.650 66.000 195.950 ;
        RECT 69.450 195.200 69.750 195.500 ;
        RECT 73.300 195.000 73.600 195.300 ;
      LAYER met3 ;
        RECT 27.100 223.850 147.200 224.350 ;
        RECT 30.600 222.950 147.200 223.450 ;
        RECT 30.600 222.050 147.200 222.550 ;
        RECT 30.600 221.150 147.200 221.650 ;
        RECT 30.600 220.250 147.200 220.750 ;
        RECT 4.000 219.350 27.600 219.850 ;
        RECT 30.600 219.350 147.200 219.850 ;
        RECT 30.600 218.450 147.200 218.950 ;
        RECT 30.600 217.550 147.200 218.050 ;
        RECT 30.600 216.700 147.200 217.150 ;
        RECT 30.600 216.650 143.850 216.700 ;
        RECT 30.600 215.750 147.200 216.250 ;
        RECT 30.600 214.850 147.200 215.350 ;
        RECT 30.600 213.950 147.200 214.450 ;
        RECT 30.600 213.050 147.200 213.550 ;
        RECT 30.600 212.150 147.200 212.650 ;
        RECT 62.650 211.750 63.150 211.800 ;
        RECT 83.000 211.750 83.500 211.800 ;
        RECT 30.600 211.350 147.200 211.750 ;
        RECT 62.650 211.300 63.150 211.350 ;
        RECT 83.000 211.300 83.500 211.350 ;
        RECT 59.150 210.950 59.650 211.000 ;
        RECT 113.400 210.950 113.900 211.000 ;
        RECT 30.600 210.550 147.200 210.950 ;
        RECT 59.150 210.500 59.650 210.550 ;
        RECT 113.400 210.500 113.900 210.550 ;
        RECT 58.250 210.150 58.750 210.200 ;
        RECT 116.150 210.150 116.650 210.200 ;
        RECT 30.600 209.750 147.200 210.150 ;
        RECT 58.250 209.700 58.750 209.750 ;
        RECT 116.150 209.700 116.650 209.750 ;
        RECT 54.550 209.350 55.050 209.400 ;
        RECT 85.800 209.350 86.300 209.400 ;
        RECT 30.600 208.950 147.200 209.350 ;
        RECT 54.550 208.900 55.050 208.950 ;
        RECT 85.800 208.900 86.300 208.950 ;
        RECT 51.550 208.550 52.050 208.600 ;
        RECT 118.900 208.550 119.400 208.600 ;
        RECT 30.600 208.150 147.200 208.550 ;
        RECT 51.550 208.100 52.050 208.150 ;
        RECT 118.900 208.100 119.400 208.150 ;
        RECT 50.550 207.750 51.050 207.800 ;
        RECT 121.650 207.750 122.150 207.800 ;
        RECT 30.600 207.350 147.200 207.750 ;
        RECT 50.550 207.300 51.050 207.350 ;
        RECT 121.650 207.300 122.150 207.350 ;
        RECT 34.850 206.950 35.350 207.000 ;
        RECT 30.600 206.550 147.200 206.950 ;
        RECT 34.850 206.500 35.350 206.550 ;
        RECT 31.700 206.150 32.200 206.200 ;
        RECT 135.400 206.150 135.900 206.200 ;
        RECT 30.600 205.750 147.200 206.150 ;
        RECT 31.700 205.700 32.200 205.750 ;
        RECT 135.400 205.700 135.900 205.750 ;
        RECT 30.800 205.350 31.300 205.400 ;
        RECT 138.200 205.350 138.700 205.400 ;
        RECT 30.600 204.950 147.200 205.350 ;
        RECT 30.800 204.900 31.300 204.950 ;
        RECT 138.200 204.900 138.700 204.950 ;
        RECT 1.000 203.800 30.500 204.300 ;
        RECT 30.800 203.150 34.800 203.650 ;
        RECT 36.750 203.150 41.050 203.650 ;
        RECT 44.150 203.500 48.500 204.000 ;
        RECT 50.550 203.500 51.500 203.600 ;
        RECT 35.950 202.600 36.450 203.100 ;
        RECT 42.100 202.650 42.600 203.150 ;
        RECT 46.000 202.250 46.500 202.750 ;
        RECT 49.650 202.650 50.150 203.150 ;
        RECT 50.550 203.100 54.900 203.500 ;
        RECT 58.250 203.250 62.560 203.750 ;
        RECT 64.700 203.200 69.000 203.700 ;
        RECT 72.250 203.450 76.650 203.900 ;
        RECT 72.250 203.400 74.000 203.450 ;
        RECT 74.550 203.400 76.650 203.450 ;
        RECT 56.100 202.700 56.600 203.200 ;
        RECT 60.100 202.550 60.950 202.950 ;
        RECT 63.650 202.700 64.150 203.200 ;
        RECT 60.450 202.450 60.950 202.550 ;
        RECT 66.650 202.250 69.050 202.650 ;
        RECT 70.250 202.600 70.750 203.100 ;
        RECT 77.950 202.650 78.450 203.150 ;
        RECT 31.700 201.750 34.200 202.250 ;
        RECT 37.750 201.700 41.500 202.200 ;
        RECT 68.550 202.150 69.050 202.250 ;
        RECT 45.000 201.450 47.600 201.950 ;
        RECT 51.550 201.550 55.450 202.050 ;
        RECT 59.150 201.500 63.050 202.000 ;
        RECT 65.700 201.450 68.250 201.950 ;
        RECT 73.250 201.600 77.400 202.100 ;
        RECT 31.700 201.050 33.000 201.450 ;
        RECT 31.700 200.950 32.200 201.050 ;
        RECT 37.900 200.700 39.250 201.100 ;
        RECT 51.650 200.850 53.000 201.250 ;
        RECT 75.900 201.200 76.400 201.300 ;
        RECT 77.000 201.200 77.500 201.300 ;
        RECT 58.200 200.600 67.950 201.000 ;
        RECT 72.350 200.800 77.500 201.200 ;
        RECT 67.450 200.500 67.950 200.600 ;
        RECT 30.900 199.950 39.950 200.350 ;
        RECT 30.900 199.900 31.300 199.950 ;
        RECT 39.450 199.850 39.950 199.950 ;
        RECT 44.900 200.150 45.400 200.250 ;
        RECT 45.950 200.150 46.450 200.250 ;
        RECT 44.900 199.750 46.450 200.150 ;
        RECT 50.700 199.900 60.200 200.300 ;
        RECT 68.500 200.150 69.000 200.250 ;
        RECT 65.750 199.750 69.000 200.150 ;
        RECT 73.400 200.050 74.700 200.450 ;
        RECT 77.900 199.750 78.400 199.850 ;
        RECT 42.000 199.400 42.500 199.500 ;
        RECT 33.050 198.850 33.550 199.400 ;
        RECT 39.200 199.000 42.500 199.400 ;
        RECT 46.400 199.400 46.900 199.450 ;
        RECT 49.600 199.400 50.100 199.500 ;
        RECT 56.050 199.400 56.550 199.500 ;
        RECT 63.650 199.400 64.150 199.500 ;
        RECT 70.200 199.405 70.700 199.500 ;
        RECT 68.100 199.400 70.700 199.405 ;
        RECT 46.400 199.000 50.100 199.400 ;
        RECT 53.000 199.000 56.550 199.400 ;
        RECT 60.500 199.000 64.150 199.400 ;
        RECT 67.100 199.000 70.700 199.400 ;
        RECT 74.700 199.350 78.400 199.750 ;
        RECT 46.400 198.950 46.900 199.000 ;
        RECT 74.150 198.650 74.550 198.850 ;
        RECT 35.900 198.550 36.400 198.650 ;
        RECT 45.900 198.600 46.400 198.650 ;
        RECT 32.700 198.150 36.400 198.550 ;
        RECT 36.900 198.200 46.400 198.600 ;
        RECT 64.700 198.250 74.550 198.650 ;
        RECT 35.900 198.100 36.400 198.150 ;
        RECT 44.050 197.450 52.850 197.850 ;
        RECT 58.500 197.700 60.200 198.100 ;
        RECT 60.400 197.050 60.900 197.150 ;
        RECT 33.050 196.650 33.550 196.750 ;
        RECT 31.100 196.250 33.550 196.650 ;
        RECT 34.850 196.550 35.350 197.050 ;
        RECT 49.600 196.900 50.100 196.950 ;
        RECT 34.900 196.400 35.300 196.550 ;
        RECT 40.900 196.400 41.400 196.900 ;
        RECT 44.400 196.500 50.100 196.900 ;
        RECT 44.400 196.400 44.900 196.500 ;
        RECT 54.600 196.450 55.000 196.700 ;
        RECT 59.150 196.650 60.900 197.050 ;
        RECT 62.600 196.450 63.100 196.950 ;
        RECT 70.150 196.850 70.650 196.950 ;
        RECT 65.050 196.450 70.650 196.850 ;
        RECT 37.750 196.000 38.250 196.050 ;
        RECT 39.450 196.000 39.950 196.100 ;
        RECT 35.900 195.800 36.400 195.900 ;
        RECT 31.700 195.400 36.400 195.800 ;
        RECT 37.750 195.600 39.950 196.000 ;
        RECT 44.950 196.050 45.450 196.100 ;
        RECT 45.850 196.050 46.350 196.150 ;
        RECT 44.950 195.650 46.350 196.050 ;
        RECT 44.950 195.600 45.450 195.650 ;
        RECT 48.800 195.600 49.300 196.100 ;
        RECT 54.550 195.950 55.050 196.450 ;
        RECT 63.650 196.050 64.150 196.150 ;
        RECT 59.150 195.650 64.150 196.050 ;
        RECT 67.450 196.000 67.950 196.100 ;
        RECT 75.900 196.000 76.400 196.500 ;
        RECT 65.650 195.600 67.950 196.000 ;
        RECT 37.750 195.550 38.250 195.600 ;
        RECT 37.250 195.150 37.650 195.250 ;
        RECT 41.850 195.150 42.450 195.350 ;
        RECT 48.850 195.250 49.250 195.600 ;
        RECT 50.850 195.250 51.350 195.300 ;
        RECT 56.050 195.250 56.550 195.350 ;
        RECT 4.000 194.400 31.200 194.900 ;
        RECT 37.250 194.850 42.450 195.150 ;
        RECT 50.850 194.850 56.550 195.250 ;
        RECT 69.300 195.150 69.800 195.650 ;
        RECT 77.850 195.350 78.350 195.450 ;
        RECT 73.250 194.950 78.350 195.350 ;
        RECT 37.250 194.650 37.750 194.850 ;
        RECT 50.850 194.800 51.350 194.850 ;
      LAYER via3 ;
        RECT 27.150 223.900 27.550 224.300 ;
        RECT 30.650 223.900 31.050 224.300 ;
        RECT 32.600 223.900 33.000 224.300 ;
        RECT 33.400 223.900 33.800 224.300 ;
        RECT 36.150 223.900 36.550 224.300 ;
        RECT 38.900 223.900 39.300 224.300 ;
        RECT 41.650 223.900 42.050 224.300 ;
        RECT 44.400 223.900 44.800 224.300 ;
        RECT 47.150 223.900 47.550 224.300 ;
        RECT 49.900 223.900 50.300 224.300 ;
        RECT 52.700 223.900 53.100 224.300 ;
        RECT 55.450 223.900 55.850 224.300 ;
        RECT 58.200 223.900 58.600 224.300 ;
        RECT 61.000 223.900 61.400 224.300 ;
        RECT 63.750 223.900 64.150 224.300 ;
        RECT 66.500 223.900 66.900 224.300 ;
        RECT 69.250 223.900 69.650 224.300 ;
        RECT 72.050 223.900 72.450 224.300 ;
        RECT 48.850 223.000 49.250 223.400 ;
        RECT 88.600 223.000 89.000 223.400 ;
        RECT 45.050 222.100 45.450 222.500 ;
        RECT 124.450 222.100 124.850 222.500 ;
        RECT 44.200 221.200 44.600 221.600 ;
        RECT 127.250 221.200 127.650 221.600 ;
        RECT 41.000 220.300 41.400 220.700 ;
        RECT 91.350 220.300 91.750 220.700 ;
        RECT 4.050 219.400 4.450 219.800 ;
        RECT 4.700 219.400 5.100 219.800 ;
        RECT 5.350 219.400 5.750 219.800 ;
        RECT 27.150 219.400 27.550 219.800 ;
        RECT 37.800 219.400 38.200 219.800 ;
        RECT 130.000 219.400 130.400 219.800 ;
        RECT 36.800 218.500 37.200 218.900 ;
        RECT 132.750 218.500 133.150 218.900 ;
        RECT 74.800 217.600 75.200 218.000 ;
        RECT 77.100 217.600 77.500 218.000 ;
        RECT 76.000 216.700 76.400 217.100 ;
        RECT 78.750 216.700 79.150 217.100 ;
        RECT 73.250 215.800 73.650 216.200 ;
        RECT 102.400 215.800 102.800 216.200 ;
        RECT 72.300 214.900 72.700 215.300 ;
        RECT 105.150 214.900 105.550 215.300 ;
        RECT 69.400 214.000 69.800 214.400 ;
        RECT 80.250 214.000 80.650 214.400 ;
        RECT 65.750 213.100 66.150 213.500 ;
        RECT 107.900 213.100 108.300 213.500 ;
        RECT 64.750 212.200 65.150 212.600 ;
        RECT 110.650 212.200 111.050 212.600 ;
        RECT 62.700 211.350 63.100 211.750 ;
        RECT 83.050 211.350 83.450 211.750 ;
        RECT 59.200 210.550 59.600 210.950 ;
        RECT 113.450 210.550 113.850 210.950 ;
        RECT 58.300 209.750 58.700 210.150 ;
        RECT 116.200 209.750 116.600 210.150 ;
        RECT 54.600 208.950 55.000 209.350 ;
        RECT 85.850 208.950 86.250 209.350 ;
        RECT 51.600 208.150 52.000 208.550 ;
        RECT 118.950 208.150 119.350 208.550 ;
        RECT 50.600 207.350 51.000 207.750 ;
        RECT 121.700 207.350 122.100 207.750 ;
        RECT 34.900 206.550 35.300 206.950 ;
        RECT 94.100 206.550 94.500 206.950 ;
        RECT 31.750 205.750 32.150 206.150 ;
        RECT 135.450 205.750 135.850 206.150 ;
        RECT 30.850 204.950 31.250 205.350 ;
        RECT 138.250 204.950 138.650 205.350 ;
        RECT 1.100 203.850 1.500 204.250 ;
        RECT 1.750 203.850 2.150 204.250 ;
        RECT 2.400 203.850 2.800 204.250 ;
        RECT 30.850 203.200 31.260 203.600 ;
        RECT 36.800 203.200 37.200 203.600 ;
        RECT 44.200 203.550 44.600 203.950 ;
        RECT 50.600 203.150 51.000 203.550 ;
        RECT 58.300 203.300 58.700 203.700 ;
        RECT 64.750 203.250 65.150 203.650 ;
        RECT 72.300 203.450 72.700 203.850 ;
        RECT 36.000 202.650 36.400 203.050 ;
        RECT 42.150 202.700 42.550 203.100 ;
        RECT 46.050 202.300 46.450 202.700 ;
        RECT 49.700 202.700 50.100 203.100 ;
        RECT 56.150 202.750 56.550 203.150 ;
        RECT 60.500 202.500 60.900 202.900 ;
        RECT 63.700 202.700 64.100 203.150 ;
        RECT 70.300 202.650 70.700 203.050 ;
        RECT 78.000 202.700 78.400 203.100 ;
        RECT 68.600 202.200 69.000 202.600 ;
        RECT 31.750 201.800 32.100 202.200 ;
        RECT 37.800 201.750 38.200 202.150 ;
        RECT 45.050 201.500 45.450 201.900 ;
        RECT 51.600 201.600 52.000 202.000 ;
        RECT 59.200 201.550 59.600 201.950 ;
        RECT 65.750 201.500 66.150 201.900 ;
        RECT 73.250 201.650 73.650 202.050 ;
        RECT 67.500 200.550 67.900 200.950 ;
        RECT 77.050 200.850 77.450 201.250 ;
        RECT 39.500 199.900 39.900 200.300 ;
        RECT 46.000 199.800 46.400 200.200 ;
        RECT 68.550 199.800 68.950 200.200 ;
        RECT 33.100 198.950 33.500 199.350 ;
        RECT 42.050 199.050 42.450 199.450 ;
        RECT 49.650 199.050 50.050 199.450 ;
        RECT 56.100 199.050 56.500 199.450 ;
        RECT 63.700 199.050 64.100 199.450 ;
        RECT 70.250 199.050 70.650 199.450 ;
        RECT 77.950 199.400 78.350 199.800 ;
        RECT 35.950 198.150 36.350 198.550 ;
        RECT 45.950 198.250 46.350 198.600 ;
        RECT 33.100 196.300 33.500 196.700 ;
        RECT 34.900 196.600 35.300 197.000 ;
        RECT 40.950 196.450 41.350 196.850 ;
        RECT 49.650 196.550 50.050 196.900 ;
        RECT 60.450 196.700 60.850 197.100 ;
        RECT 62.650 196.500 63.050 196.900 ;
        RECT 70.200 196.500 70.600 196.900 ;
        RECT 35.950 195.450 36.350 195.850 ;
        RECT 37.800 195.600 38.200 196.000 ;
        RECT 39.500 195.650 39.900 196.050 ;
        RECT 45.900 195.700 46.300 196.100 ;
        RECT 48.850 195.650 49.250 196.050 ;
        RECT 54.600 196.000 55.000 196.400 ;
        RECT 63.700 195.700 64.100 196.100 ;
        RECT 67.500 195.650 67.900 196.050 ;
        RECT 75.950 196.050 76.350 196.450 ;
        RECT 42.000 194.900 42.400 195.300 ;
        RECT 4.100 194.450 4.500 194.850 ;
        RECT 4.750 194.450 5.150 194.850 ;
        RECT 5.400 194.450 5.800 194.850 ;
        RECT 56.100 194.900 56.500 195.300 ;
        RECT 69.350 195.200 69.750 195.600 ;
        RECT 77.900 195.000 78.300 195.400 ;
      LAYER met4 ;
        RECT 30.650 224.760 30.670 224.850 ;
        RECT 30.970 224.760 31.050 224.850 ;
        RECT 30.650 224.350 31.050 224.760 ;
        RECT 33.400 224.760 33.430 224.850 ;
        RECT 33.730 224.760 33.800 224.850 ;
        RECT 33.400 224.350 33.800 224.760 ;
        RECT 36.150 224.760 36.190 224.850 ;
        RECT 36.490 224.760 36.550 224.850 ;
        RECT 36.150 224.350 36.550 224.760 ;
        RECT 38.900 224.760 38.950 224.850 ;
        RECT 39.250 224.760 39.300 224.850 ;
        RECT 38.900 224.350 39.300 224.760 ;
        RECT 41.650 224.760 41.710 224.850 ;
        RECT 42.010 224.760 42.050 224.850 ;
        RECT 41.650 224.350 42.050 224.760 ;
        RECT 44.400 224.760 44.470 224.850 ;
        RECT 44.770 224.760 44.800 224.850 ;
        RECT 44.400 224.350 44.800 224.760 ;
        RECT 47.150 224.760 47.230 224.850 ;
        RECT 47.530 224.760 47.550 224.850 ;
        RECT 47.150 224.350 47.550 224.760 ;
        RECT 49.900 224.760 49.990 224.850 ;
        RECT 50.290 224.760 50.300 224.850 ;
        RECT 49.900 224.350 50.300 224.760 ;
        RECT 52.700 224.760 52.750 224.950 ;
        RECT 53.050 224.760 53.100 224.950 ;
        RECT 52.700 224.350 53.100 224.760 ;
        RECT 55.450 224.760 55.510 224.900 ;
        RECT 55.810 224.760 55.850 224.900 ;
        RECT 55.450 224.350 55.850 224.760 ;
        RECT 58.200 224.760 58.270 224.900 ;
        RECT 58.570 224.760 58.600 224.900 ;
        RECT 58.200 224.350 58.600 224.760 ;
        RECT 61.000 224.760 61.030 224.900 ;
        RECT 61.330 224.760 61.400 224.900 ;
        RECT 61.000 224.350 61.400 224.760 ;
        RECT 63.750 224.760 63.790 224.950 ;
        RECT 64.090 224.760 64.150 224.950 ;
        RECT 63.750 224.350 64.150 224.760 ;
        RECT 66.500 224.760 66.550 224.900 ;
        RECT 66.850 224.760 66.900 224.900 ;
        RECT 66.500 224.350 66.900 224.760 ;
        RECT 69.250 224.760 69.310 225.050 ;
        RECT 69.610 224.760 69.650 225.050 ;
        RECT 69.250 224.350 69.650 224.760 ;
        RECT 72.050 224.760 72.070 224.900 ;
        RECT 72.370 224.760 72.450 224.900 ;
        RECT 72.050 224.350 72.450 224.760 ;
        RECT 74.800 224.760 74.830 224.900 ;
        RECT 75.130 224.760 75.200 224.900 ;
        RECT 27.100 223.850 27.600 224.350 ;
        RECT 30.600 223.850 31.100 224.350 ;
        RECT 32.550 223.850 33.050 224.350 ;
        RECT 33.350 223.850 33.850 224.350 ;
        RECT 36.100 223.850 36.600 224.350 ;
        RECT 38.850 223.850 39.350 224.350 ;
        RECT 41.600 223.850 42.100 224.350 ;
        RECT 44.350 223.850 44.850 224.350 ;
        RECT 47.100 223.850 47.600 224.350 ;
        RECT 49.850 223.850 50.350 224.350 ;
        RECT 52.650 223.850 53.150 224.350 ;
        RECT 55.400 223.850 55.900 224.350 ;
        RECT 58.150 223.850 58.650 224.350 ;
        RECT 60.950 223.850 61.450 224.350 ;
        RECT 63.700 223.850 64.200 224.350 ;
        RECT 66.450 223.850 66.950 224.350 ;
        RECT 69.200 223.850 69.700 224.350 ;
        RECT 72.000 223.850 72.500 224.350 ;
        RECT 27.150 219.850 27.550 223.850 ;
        RECT 27.100 219.350 27.600 219.850 ;
        RECT 31.700 205.700 32.200 206.200 ;
        RECT 30.800 204.900 31.300 205.400 ;
        RECT 30.850 203.650 31.250 204.900 ;
        RECT 30.800 203.150 31.300 203.650 ;
        RECT 31.750 202.250 32.150 205.700 ;
        RECT 32.600 204.750 33.000 223.850 ;
        RECT 48.800 222.950 49.300 223.450 ;
        RECT 45.000 222.050 45.500 222.550 ;
        RECT 44.150 221.150 44.650 221.650 ;
        RECT 40.950 220.250 41.450 220.750 ;
        RECT 37.750 219.350 38.250 219.850 ;
        RECT 36.750 218.450 37.250 218.950 ;
        RECT 34.850 206.500 35.350 207.000 ;
        RECT 32.600 204.450 33.500 204.750 ;
        RECT 31.700 201.750 32.150 202.250 ;
        RECT 33.050 199.400 33.500 204.450 ;
        RECT 33.050 198.850 33.550 199.400 ;
        RECT 33.150 196.750 33.550 198.850 ;
        RECT 34.900 197.050 35.300 206.500 ;
        RECT 36.800 203.650 37.200 218.450 ;
        RECT 36.750 203.150 37.250 203.650 ;
        RECT 35.950 202.600 36.450 203.100 ;
        RECT 36.000 198.650 36.400 202.600 ;
        RECT 37.800 202.200 38.200 219.350 ;
        RECT 37.750 201.700 38.250 202.200 ;
        RECT 39.450 199.850 39.950 200.350 ;
        RECT 35.900 198.100 36.400 198.650 ;
        RECT 33.050 196.250 33.550 196.750 ;
        RECT 34.850 196.550 35.350 197.050 ;
        RECT 36.000 196.250 36.400 198.100 ;
        RECT 35.450 195.600 36.400 196.250 ;
        RECT 39.550 196.100 39.950 199.850 ;
        RECT 41.000 196.900 41.400 220.250 ;
        RECT 44.200 204.000 44.600 221.150 ;
        RECT 44.150 203.500 44.650 204.000 ;
        RECT 42.100 202.650 42.600 203.150 ;
        RECT 42.200 199.500 42.500 202.650 ;
        RECT 45.050 201.950 45.450 222.050 ;
        RECT 46.000 202.250 46.500 202.750 ;
        RECT 45.000 201.450 45.600 201.950 ;
        RECT 46.050 200.250 46.450 202.250 ;
        RECT 45.950 199.750 46.450 200.250 ;
        RECT 42.000 199.000 42.500 199.500 ;
        RECT 40.900 196.400 41.400 196.900 ;
        RECT 35.900 195.400 36.400 195.600 ;
        RECT 37.750 195.550 38.250 196.050 ;
        RECT 39.450 195.600 39.950 196.100 ;
        RECT 42.050 195.350 42.450 199.000 ;
        RECT 45.900 198.200 46.400 198.650 ;
        RECT 45.950 196.150 46.350 198.200 ;
        RECT 45.850 195.650 46.350 196.150 ;
        RECT 48.850 196.100 49.250 222.950 ;
        RECT 74.800 218.050 75.200 224.760 ;
        RECT 77.550 224.760 77.590 224.900 ;
        RECT 77.890 224.760 77.950 224.900 ;
        RECT 77.550 224.350 77.950 224.760 ;
        RECT 80.250 224.760 80.350 225.500 ;
        RECT 83.050 224.760 83.110 224.950 ;
        RECT 83.410 224.760 83.450 224.950 ;
        RECT 77.550 223.850 79.150 224.350 ;
        RECT 74.750 217.550 75.250 218.050 ;
        RECT 77.050 217.550 77.550 218.050 ;
        RECT 75.950 216.650 76.450 217.150 ;
        RECT 73.200 215.750 73.700 216.250 ;
        RECT 72.250 214.850 72.750 215.350 ;
        RECT 69.350 213.950 69.850 214.450 ;
        RECT 65.700 213.050 66.200 213.550 ;
        RECT 64.700 212.150 65.200 212.650 ;
        RECT 62.650 211.300 63.150 211.800 ;
        RECT 59.150 210.500 59.650 211.000 ;
        RECT 58.250 209.700 58.750 210.200 ;
        RECT 54.550 208.900 55.050 209.400 ;
        RECT 51.550 208.100 52.050 208.600 ;
        RECT 50.550 207.300 51.050 207.800 ;
        RECT 50.600 203.600 51.000 207.300 ;
        RECT 49.650 202.650 50.150 203.150 ;
        RECT 50.550 203.100 51.100 203.600 ;
        RECT 49.700 199.500 50.100 202.650 ;
        RECT 51.600 202.050 52.000 208.100 ;
        RECT 51.550 201.550 52.050 202.050 ;
        RECT 49.600 199.000 50.100 199.500 ;
        RECT 49.700 196.950 50.100 199.000 ;
        RECT 49.600 196.500 50.100 196.950 ;
        RECT 54.600 196.450 55.000 208.900 ;
        RECT 58.300 203.750 58.700 209.700 ;
        RECT 58.250 203.250 58.850 203.750 ;
        RECT 56.100 202.700 56.600 203.200 ;
        RECT 56.150 199.500 56.550 202.700 ;
        RECT 59.200 202.000 59.600 210.500 ;
        RECT 60.450 202.450 60.950 202.950 ;
        RECT 59.150 201.500 59.700 202.000 ;
        RECT 56.050 199.000 56.550 199.500 ;
        RECT 48.800 195.600 49.300 196.100 ;
        RECT 54.550 195.950 55.050 196.450 ;
        RECT 56.150 195.350 56.550 199.000 ;
        RECT 60.500 197.150 60.900 202.450 ;
        RECT 60.400 196.650 60.900 197.150 ;
        RECT 62.700 196.950 63.100 211.300 ;
        RECT 64.750 203.700 65.150 212.150 ;
        RECT 64.700 203.200 65.250 203.700 ;
        RECT 63.650 202.650 64.150 203.200 ;
        RECT 63.750 199.500 64.150 202.650 ;
        RECT 65.750 201.950 66.150 213.050 ;
        RECT 68.550 202.150 69.050 202.650 ;
        RECT 65.700 201.450 66.245 201.950 ;
        RECT 67.450 200.500 67.950 201.000 ;
        RECT 63.650 199.000 64.150 199.500 ;
        RECT 62.600 196.450 63.100 196.950 ;
        RECT 63.750 196.150 64.150 199.000 ;
        RECT 63.650 195.650 64.150 196.150 ;
        RECT 67.550 196.100 67.950 200.500 ;
        RECT 68.600 200.250 69.000 202.150 ;
        RECT 68.500 199.750 69.000 200.250 ;
        RECT 67.450 195.600 67.950 196.100 ;
        RECT 69.400 195.650 69.800 213.950 ;
        RECT 72.300 203.900 72.700 214.850 ;
        RECT 72.250 203.400 72.950 203.900 ;
        RECT 70.250 202.600 70.750 203.100 ;
        RECT 70.300 199.500 70.700 202.600 ;
        RECT 73.250 202.250 73.650 215.750 ;
        RECT 73.200 201.600 73.700 202.250 ;
        RECT 76.000 201.300 76.400 216.650 ;
        RECT 77.100 201.300 77.500 217.550 ;
        RECT 78.750 217.150 79.150 223.850 ;
        RECT 78.700 216.650 79.200 217.150 ;
        RECT 80.250 214.450 80.650 224.760 ;
        RECT 80.200 213.950 80.700 214.450 ;
        RECT 83.050 211.800 83.450 224.760 ;
        RECT 85.850 224.760 85.870 224.900 ;
        RECT 86.170 224.760 86.250 224.900 ;
        RECT 83.000 211.300 83.500 211.800 ;
        RECT 85.850 209.400 86.250 224.760 ;
        RECT 88.600 224.760 88.630 224.900 ;
        RECT 88.930 224.760 89.000 224.900 ;
        RECT 88.600 223.450 89.000 224.760 ;
        RECT 91.350 224.760 91.390 224.900 ;
        RECT 91.690 224.760 91.750 224.900 ;
        RECT 88.550 222.950 89.050 223.450 ;
        RECT 91.350 220.750 91.750 224.760 ;
        RECT 94.100 224.760 94.150 224.900 ;
        RECT 94.450 224.760 94.500 224.900 ;
        RECT 91.300 220.250 91.800 220.750 ;
        RECT 85.800 208.900 86.300 209.400 ;
        RECT 94.100 207.000 94.500 224.760 ;
        RECT 102.400 224.760 102.430 224.900 ;
        RECT 102.730 224.760 102.800 224.900 ;
        RECT 102.400 216.250 102.800 224.760 ;
        RECT 105.150 224.760 105.190 224.850 ;
        RECT 105.490 224.760 105.550 224.850 ;
        RECT 102.350 215.750 102.850 216.250 ;
        RECT 105.150 215.350 105.550 224.760 ;
        RECT 107.900 224.760 107.950 224.900 ;
        RECT 108.250 224.760 108.300 224.900 ;
        RECT 105.100 214.850 105.600 215.350 ;
        RECT 107.900 213.550 108.300 224.760 ;
        RECT 110.650 224.760 110.710 224.850 ;
        RECT 111.010 224.760 111.050 224.850 ;
        RECT 107.850 213.050 108.350 213.550 ;
        RECT 110.650 212.650 111.050 224.760 ;
        RECT 113.450 224.760 113.470 224.900 ;
        RECT 113.770 224.760 113.850 224.900 ;
        RECT 110.600 212.150 111.100 212.650 ;
        RECT 113.450 211.000 113.850 224.760 ;
        RECT 116.200 224.760 116.230 224.850 ;
        RECT 116.530 224.760 116.600 224.850 ;
        RECT 113.400 210.500 113.900 211.000 ;
        RECT 116.200 210.200 116.600 224.760 ;
        RECT 118.950 224.760 118.990 224.900 ;
        RECT 119.290 224.760 119.350 224.900 ;
        RECT 116.150 209.700 116.650 210.200 ;
        RECT 118.950 208.600 119.350 224.760 ;
        RECT 121.700 224.760 121.750 224.900 ;
        RECT 122.050 224.760 122.100 224.900 ;
        RECT 118.900 208.100 119.400 208.600 ;
        RECT 121.700 207.800 122.100 224.760 ;
        RECT 124.450 224.760 124.510 224.900 ;
        RECT 124.810 224.760 124.850 224.900 ;
        RECT 124.450 222.550 124.850 224.760 ;
        RECT 127.250 224.760 127.270 224.900 ;
        RECT 127.570 224.760 127.650 224.900 ;
        RECT 124.400 222.050 124.900 222.550 ;
        RECT 127.250 221.650 127.650 224.760 ;
        RECT 130.000 224.760 130.030 224.850 ;
        RECT 130.330 224.760 130.400 224.850 ;
        RECT 127.200 221.150 127.700 221.650 ;
        RECT 130.000 219.850 130.400 224.760 ;
        RECT 132.750 224.760 132.790 224.850 ;
        RECT 133.090 224.760 133.150 224.850 ;
        RECT 129.950 219.350 130.450 219.850 ;
        RECT 132.750 218.950 133.150 224.760 ;
        RECT 135.450 224.760 135.550 225.300 ;
        RECT 138.250 224.760 138.310 224.900 ;
        RECT 138.610 224.760 138.650 224.900 ;
        RECT 132.700 218.450 133.200 218.950 ;
        RECT 121.650 207.300 122.150 207.800 ;
        RECT 94.050 206.500 94.550 207.000 ;
        RECT 135.450 206.200 135.850 224.760 ;
        RECT 135.400 205.700 135.900 206.200 ;
        RECT 138.250 205.400 138.650 224.760 ;
        RECT 138.200 204.900 138.700 205.400 ;
        RECT 77.950 202.650 78.450 203.150 ;
        RECT 75.900 200.800 76.400 201.300 ;
        RECT 77.000 200.800 77.500 201.300 ;
        RECT 70.200 199.000 70.700 199.500 ;
        RECT 70.250 196.950 70.650 199.000 ;
        RECT 70.150 196.450 70.650 196.950 ;
        RECT 76.000 196.500 76.400 200.800 ;
        RECT 78.000 199.850 78.400 202.650 ;
        RECT 77.900 199.350 78.400 199.850 ;
        RECT 75.900 196.000 76.400 196.500 ;
        RECT 41.850 194.850 42.450 195.350 ;
        RECT 56.050 194.850 56.550 195.350 ;
        RECT 69.300 195.150 69.800 195.650 ;
        RECT 77.950 195.450 78.350 199.350 ;
        RECT 77.850 194.950 78.350 195.450 ;
  END
END tt_um_carry_ripple_7_bit
END LIBRARY

