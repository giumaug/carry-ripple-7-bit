magic
tech sky130A
magscale 1 2
timestamp 1740396551
<< nwell >>
rect -40 260 9580 592
rect 2540 -100 2710 -78
rect 2540 -400 2630 -100
rect 2540 -420 2710 -400
rect 3234 -409 3270 -88
rect 3870 -409 3937 -88
rect 4543 -409 4568 -88
rect 5185 -406 5245 -88
rect 5394 -398 5460 -86
rect 5394 -406 5580 -398
rect 5185 -407 5580 -406
rect 6045 -407 6090 -86
rect 6700 -407 6754 -86
rect 7365 -407 7395 -86
rect 8013 -407 8068 -86
rect 8200 -90 8370 -80
rect 8200 -400 8300 -90
rect 5188 -410 5580 -407
rect 8200 -410 8370 -400
rect 8895 -407 8952 -86
rect 5400 -760 5570 -750
rect 671 -1081 692 -760
rect 1120 -1081 1182 -760
rect 1880 -1081 1940 -760
rect 2360 -1081 2417 -760
rect 2570 -1080 2630 -760
rect 5400 -1080 5450 -760
rect 2570 -1090 2750 -1080
rect 5400 -1090 5570 -1080
rect 6155 -1081 6184 -760
rect 7460 -1081 7484 -760
rect 8224 -1081 8276 -760
rect 8986 -1081 9131 -760
<< pwell >>
rect 1109 -49 1235 60
rect 1665 -48 1720 48
<< locali >>
rect 454 527 502 561
rect 1121 527 1217 561
rect 1665 527 1719 561
rect 2349 527 2453 561
rect 2532 527 2668 561
rect 3115 527 3233 561
rect 3866 527 3973 561
rect 4427 527 4530 561
rect 5170 527 5282 561
rect 5363 527 5481 561
rect 5928 527 6044 561
rect 6675 527 6792 561
rect 7246 527 7352 561
rect 7990 527 8104 561
rect 8184 527 8313 561
rect 8759 527 8894 561
rect 10 280 90 300
rect 10 240 30 280
rect 70 240 90 280
rect 10 220 90 240
rect 2026 249 2101 260
rect 2026 243 2051 249
rect 2085 243 2101 249
rect 437 -17 504 17
rect 1117 -17 1221 17
rect 1656 -18 1720 17
rect 2348 -17 2457 17
rect 2526 -17 2661 17
rect 3115 -17 3235 17
rect 3863 -17 3973 17
rect 4417 -17 4534 17
rect 5170 -17 5285 17
rect 5359 -17 5483 17
rect 5925 -17 6047 17
rect 6678 -17 6794 17
rect 7237 -17 7354 17
rect 7981 -17 8104 17
rect 8178 -17 8315 17
rect 8768 -17 8894 17
rect 5110 -109 5280 -104
rect 529 -145 624 -111
rect 1169 -145 1231 -109
rect 1756 -143 1842 -109
rect 2388 -143 2452 -109
rect 2523 -143 2664 -109
rect 3208 -143 3316 -109
rect 3828 -143 3974 -109
rect 4513 -143 4604 -109
rect 5110 -120 5282 -109
rect 5149 -141 5282 -120
rect 5367 -141 5487 -107
rect 6027 -141 6121 -107
rect 6655 -141 6799 -107
rect 7337 -141 7433 -107
rect 7977 -141 8103 -107
rect 8183 -141 8314 -107
rect 8857 -141 8987 -107
rect 545 -689 624 -655
rect 1155 -660 1220 -650
rect 5126 -653 5281 -651
rect 1163 -687 1217 -660
rect 1762 -687 1843 -653
rect 2383 -687 2453 -653
rect 2533 -687 2665 -653
rect 3200 -687 3293 -653
rect 3830 -687 3976 -653
rect 4502 -687 4603 -653
rect 5126 -686 5285 -653
rect 5362 -685 5484 -651
rect 6027 -686 6126 -651
rect 6661 -685 6793 -651
rect 7333 -685 7433 -651
rect 7974 -685 8107 -651
rect 8189 -685 8313 -651
rect 8859 -685 8997 -651
rect 5126 -687 5281 -686
rect 626 -815 732 -781
rect 1092 -815 1222 -781
rect 1844 -815 1977 -781
rect 2332 -815 2451 -781
rect 2537 -815 2660 -781
rect 3293 -815 3364 -781
rect 3895 -815 3973 -781
rect 4600 -815 4692 -781
rect 5233 -815 5283 -781
rect 5369 -815 5490 -781
rect 6111 -815 6226 -781
rect 6763 -815 6792 -781
rect 7425 -815 7523 -781
rect 8060 -815 8106 -781
rect 8187 -815 8318 -781
rect 8944 -815 9174 -781
rect 632 -1359 732 -1325
rect 1087 -1359 1224 -1325
rect 1851 -1359 1975 -1325
rect 2330 -1359 2455 -1325
rect 2528 -1359 2666 -1325
rect 3293 -1359 3363 -1325
rect 3902 -1360 3974 -1325
rect 4603 -1359 4694 -1325
rect 5228 -1359 5285 -1325
rect 5368 -1359 5484 -1325
rect 6113 -1359 6225 -1325
rect 6758 -1359 6811 -1325
rect 7426 -1359 7524 -1325
rect 8062 -1359 8110 -1325
rect 8186 -1359 8313 -1325
rect 8945 -1359 9174 -1325
<< viali >>
rect 30 240 70 280
rect 571 270 606 306
rect 210 220 250 260
rect 680 218 716 253
rect 1240 230 1280 270
rect 1429 215 1463 249
rect 1915 215 1950 251
rect 2051 215 2085 249
rect 2690 220 2730 260
rect 2873 223 2907 258
rect 3320 215 3356 250
rect 3430 210 3470 250
rect 3990 220 4030 260
rect 4720 210 4760 250
<< metal1 >>
rect 444 496 498 592
rect 1115 496 1218 592
rect 1669 496 1720 592
rect 2354 496 2456 592
rect 2537 496 2661 592
rect 3110 496 3238 592
rect 3851 496 3977 592
rect 4423 496 4532 592
rect 5167 496 5282 592
rect 5367 496 5484 592
rect 5934 496 6044 592
rect 6679 496 6791 592
rect 7240 496 7354 592
rect 7987 496 8105 592
rect 8188 496 8312 592
rect 8765 496 8898 592
rect 550 306 619 330
rect 10 290 90 300
rect 10 230 20 290
rect 80 230 90 290
rect 10 220 90 230
rect 190 260 270 290
rect 550 270 571 306
rect 606 270 619 306
rect 660 280 740 290
rect 660 270 670 280
rect 550 260 619 270
rect 190 220 210 260
rect 250 220 270 260
rect 190 210 270 220
rect 650 220 670 270
rect 730 270 740 280
rect 1200 280 1310 290
rect 730 220 760 270
rect 650 218 680 220
rect 716 218 760 220
rect 650 210 760 218
rect 1200 220 1210 280
rect 1270 270 1310 280
rect 1900 270 1980 280
rect 1280 230 1310 270
rect 1270 220 1310 230
rect 1200 210 1310 220
rect 1413 249 1490 270
rect 1413 215 1429 249
rect 1463 215 1490 249
rect 1413 190 1490 215
rect 1900 210 1910 270
rect 1970 210 1980 270
rect 2680 270 2760 280
rect 2026 250 2100 258
rect 1900 200 1980 210
rect 2020 249 2100 250
rect 2020 240 2051 249
rect 2085 240 2100 249
rect 2020 180 2030 240
rect 2090 180 2100 240
rect 2680 210 2690 270
rect 2750 210 2760 270
rect 2680 200 2760 210
rect 2850 270 2930 280
rect 3410 270 3490 280
rect 2850 210 2860 270
rect 2920 210 2930 270
rect 3313 260 3362 270
rect 2850 190 2930 210
rect 3280 250 3362 260
rect 3280 215 3320 250
rect 3356 215 3362 250
rect 3280 199 3362 215
rect 3410 210 3420 270
rect 3480 210 3490 270
rect 3410 200 3490 210
rect 3960 270 4040 280
rect 3960 210 3970 270
rect 4030 210 4040 270
rect 3960 200 4040 210
rect 4700 210 4720 270
rect 4780 210 4800 270
rect 4700 200 4800 210
rect 3280 190 3360 199
rect 2020 170 2100 180
rect 447 -49 518 48
rect 1114 -49 1223 48
rect 1665 -48 1720 48
rect 2352 17 2461 48
rect 2348 -17 2461 17
rect 2352 -49 2461 -17
rect 2535 -48 2666 48
rect 3111 -48 3238 48
rect 3867 -48 3973 48
rect 4423 -14 4532 48
rect 4422 -48 4651 -14
rect 5166 -48 5285 48
rect 5365 -48 5486 48
rect 5933 -48 6045 48
rect 6675 -48 6794 48
rect 7244 -48 7357 48
rect 7986 -48 8108 48
rect 8185 -48 8314 48
rect 8761 -48 8894 48
rect 541 -176 635 -80
rect 1154 -174 1219 -80
rect 1762 -174 1846 -78
rect 2381 -174 2454 -78
rect 2532 -174 2664 -78
rect 3200 -174 3300 -78
rect 3835 -174 3976 -78
rect 4504 -174 4606 -78
rect 5144 -172 5283 -78
rect 5361 -172 5487 -76
rect 6023 -172 6124 -76
rect 6665 -172 6794 -76
rect 7334 -172 7431 -76
rect 7974 -172 8104 -76
rect 8186 -172 8313 -76
rect 8845 -172 8988 -76
rect 537 -720 623 -624
rect 1167 -718 1217 -624
rect 1755 -718 1843 -622
rect 2386 -718 2453 -622
rect 2535 -718 2666 -622
rect 3204 -718 3295 -622
rect 3834 -718 3976 -622
rect 4515 -718 4604 -622
rect 5144 -720 5283 -620
rect 5365 -716 5487 -620
rect 6024 -716 6125 -620
rect 6666 -716 6795 -620
rect 7336 -716 7436 -620
rect 7977 -716 8107 -620
rect 8186 -716 8315 -620
rect 8856 -716 8992 -620
rect 634 -846 735 -750
rect 1086 -846 1219 -750
rect 1851 -846 1983 -750
rect 2335 -846 2454 -750
rect 2535 -846 2662 -750
rect 3298 -846 3364 -750
rect 3902 -846 3974 -750
rect 4606 -846 4693 -750
rect 5232 -846 5284 -750
rect 5366 -846 5484 -750
rect 6116 -846 6225 -750
rect 6756 -846 6806 -750
rect 7424 -846 7523 -750
rect 8065 -846 8112 -750
rect 8181 -846 8314 -750
rect 8937 -846 9175 -750
rect 637 -1390 734 -1294
rect 1090 -1390 1222 -1294
rect 1854 -1390 1980 -1294
rect 2336 -1390 2454 -1294
rect 2534 -1390 2665 -1294
rect 3297 -1390 3364 -1294
rect 3906 -1390 3978 -1294
rect 4606 -1390 4696 -1294
rect 5233 -1390 5292 -1294
rect 5364 -1390 5488 -1294
rect 6116 -1390 6226 -1294
rect 6765 -1390 6813 -1294
rect 7425 -1390 7527 -1294
rect 8065 -1390 8105 -1294
rect 8188 -1390 8316 -1294
rect 8944 -1390 9170 -1294
<< via1 >>
rect 20 280 80 290
rect 20 240 30 280
rect 30 240 70 280
rect 70 240 80 280
rect 20 230 80 240
rect 670 253 730 280
rect 670 220 680 253
rect 680 220 716 253
rect 716 220 730 253
rect 1210 270 1270 280
rect 1210 230 1240 270
rect 1240 230 1270 270
rect 1210 220 1270 230
rect 1910 251 1970 270
rect 1910 215 1915 251
rect 1915 215 1950 251
rect 1950 215 1970 251
rect 1910 210 1970 215
rect 2030 215 2051 240
rect 2051 215 2085 240
rect 2085 215 2090 240
rect 2030 180 2090 215
rect 2690 260 2750 270
rect 2690 220 2730 260
rect 2730 220 2750 260
rect 2690 210 2750 220
rect 2860 258 2920 270
rect 2860 223 2873 258
rect 2873 223 2907 258
rect 2907 223 2920 258
rect 2860 210 2920 223
rect 3420 250 3480 270
rect 3420 210 3430 250
rect 3430 210 3470 250
rect 3470 210 3480 250
rect 3970 260 4030 270
rect 3970 220 3990 260
rect 3990 220 4030 260
rect 3970 210 4030 220
rect 4720 250 4780 270
rect 4720 210 4760 250
rect 4760 210 4780 250
<< metal2 >>
rect 2680 500 2760 530
rect 0 440 100 460
rect 0 380 20 440
rect 80 380 100 440
rect 0 360 100 380
rect 660 440 740 460
rect 720 380 740 440
rect 10 290 90 360
rect 10 230 20 290
rect 80 230 90 290
rect 10 220 90 230
rect 190 180 270 290
rect 550 180 630 330
rect 660 280 740 380
rect 1190 440 1280 460
rect 1190 380 1210 440
rect 1270 380 1280 440
rect 1190 360 1280 380
rect 660 220 670 280
rect 730 220 740 280
rect 660 210 740 220
rect 1200 280 1280 360
rect 1900 430 1990 460
rect 1900 370 1910 430
rect 1970 370 1990 430
rect 1900 290 1990 370
rect 1200 220 1210 280
rect 1270 220 1280 280
rect 1890 270 1990 290
rect 1200 210 1280 220
rect 180 160 270 180
rect 180 100 190 160
rect 250 100 270 160
rect 180 80 270 100
rect 540 160 630 180
rect 1413 170 1490 270
rect 1890 210 1910 270
rect 1970 210 1990 270
rect 2680 440 2690 500
rect 2750 440 2760 500
rect 2680 270 2760 440
rect 3410 500 3490 530
rect 3410 440 3420 500
rect 3480 440 3490 500
rect 1890 190 1990 210
rect 2020 240 2100 250
rect 540 100 560 160
rect 620 100 630 160
rect 540 80 630 100
rect 1390 150 1490 170
rect 1390 90 1410 150
rect 1470 90 1490 150
rect 1390 70 1490 90
rect 2020 180 2030 240
rect 2090 180 2100 240
rect 2680 210 2690 270
rect 2750 210 2760 270
rect 2680 200 2760 210
rect 2850 270 2930 279
rect 2850 210 2860 270
rect 2920 210 2930 270
rect 3410 270 3490 440
rect 2020 141 2100 180
rect 2080 80 2100 141
rect 2020 69 2100 80
rect 2850 100 2930 210
rect 2850 40 2860 100
rect 2920 40 2930 100
rect 2850 20 2930 40
rect 3280 100 3360 260
rect 3410 210 3420 270
rect 3480 210 3490 270
rect 3410 200 3490 210
rect 3960 430 4040 450
rect 3960 370 3970 430
rect 4030 370 4040 430
rect 3960 270 4040 370
rect 4720 270 4800 320
rect 3960 210 3970 270
rect 4030 210 4040 270
rect 3960 200 4040 210
rect 4700 210 4720 270
rect 4780 210 4800 270
rect 4700 200 4800 210
rect 3280 40 3290 100
rect 3350 40 3360 100
rect 3280 20 3360 40
<< via2 >>
rect 20 380 80 440
rect 660 380 720 440
rect 1210 380 1270 440
rect 1910 370 1970 430
rect 190 100 250 160
rect 2690 440 2750 500
rect 3420 440 3480 500
rect 560 100 620 160
rect 1410 90 1470 150
rect 2020 80 2080 141
rect 2860 40 2920 100
rect 3970 370 4030 430
rect 3290 40 3350 100
<< metal3 >>
rect 2670 520 3540 530
rect 0 450 800 460
rect 0 370 10 450
rect 92 440 800 450
rect 92 380 660 440
rect 720 380 800 440
rect 92 370 800 380
rect 0 360 800 370
rect 1190 450 2050 460
rect 1190 370 1200 450
rect 1280 430 2050 450
rect 2670 440 2680 520
rect 2760 500 3540 520
rect 2760 440 3420 500
rect 3480 440 3540 500
rect 2670 430 3540 440
rect 3950 440 4140 450
rect 1280 370 1910 430
rect 1970 370 2050 430
rect 1190 360 2050 370
rect 3950 360 3960 440
rect 4040 430 4140 440
rect 4040 360 4820 430
rect 3950 350 4820 360
rect 180 170 680 180
rect 180 90 190 170
rect 260 160 680 170
rect 260 100 560 160
rect 620 100 680 160
rect 260 90 680 100
rect 180 80 680 90
rect 1390 160 2140 170
rect 1390 80 1400 160
rect 1480 141 2140 160
rect 1480 80 2020 141
rect 2080 80 2140 141
rect 1390 70 2140 80
rect 2840 110 3360 120
rect 2840 30 2850 110
rect 2930 100 3360 110
rect 2930 40 3290 100
rect 3350 40 3360 100
rect 2930 30 3360 40
rect 2840 20 3360 30
<< via3 >>
rect 10 440 92 450
rect 10 380 20 440
rect 20 380 80 440
rect 80 380 92 440
rect 10 370 92 380
rect 1200 440 1280 450
rect 1200 380 1210 440
rect 1210 380 1270 440
rect 1270 380 1280 440
rect 2680 500 2760 520
rect 2680 440 2690 500
rect 2690 440 2750 500
rect 2750 440 2760 500
rect 1200 370 1280 380
rect 3960 430 4040 440
rect 3960 370 3970 430
rect 3970 370 4030 430
rect 4030 370 4040 430
rect 3960 360 4040 370
rect 190 160 260 170
rect 190 100 250 160
rect 250 100 260 160
rect 190 90 260 100
rect 1400 150 1480 160
rect 1400 90 1410 150
rect 1410 90 1470 150
rect 1470 90 1480 150
rect 1400 80 1480 90
rect 2850 100 2930 110
rect 2850 40 2860 100
rect 2860 40 2920 100
rect 2920 40 2930 100
rect 2850 30 2930 40
<< metal4 >>
rect 10 460 90 640
rect 0 450 100 460
rect 0 370 10 450
rect 92 370 100 450
rect 0 360 100 370
rect 190 180 270 630
rect 1200 460 1280 650
rect 1190 450 1290 460
rect 1190 370 1200 450
rect 1280 370 1290 450
rect 1190 360 1290 370
rect 180 170 270 180
rect 1400 170 1480 670
rect 2680 530 2760 640
rect 2670 520 2770 530
rect 2670 440 2680 520
rect 2760 440 2770 520
rect 2670 430 2770 440
rect 180 90 190 170
rect 260 90 270 170
rect 180 80 270 90
rect 1390 160 1490 170
rect 1390 80 1400 160
rect 1480 80 1490 160
rect 2850 120 2930 640
rect 3960 450 4040 640
rect 3950 440 4060 450
rect 3950 360 3960 440
rect 4040 360 4060 440
rect 3950 350 4060 360
rect 1390 70 1490 80
rect 2840 110 2960 120
rect 2840 30 2850 110
rect 2930 30 2960 110
rect 2840 20 2960 30
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_0
timestamp 1691611044
transform 1 0 0 0 1 -672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_1
timestamp 1691611044
transform 1 0 1214 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_2
timestamp 1691611044
transform 1 0 2658 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_3
timestamp 1691611044
transform 1 0 3968 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_4
timestamp 1691611044
transform 1 0 5478 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_5
timestamp 1691611044
transform 1 0 6788 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_6
timestamp 1691611044
transform 1 0 8310 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0
timestamp 1691611044
transform 1 0 0 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_1
timestamp 1691611044
transform 1 0 1214 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_2
timestamp 1691611044
transform 1 0 2658 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_3
timestamp 1691611044
transform 1 0 3968 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_4
timestamp 1691611044
transform 1 0 5478 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_5
timestamp 1691611044
transform 1 0 6788 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_6
timestamp 1691611044
transform 1 0 8310 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0
timestamp 1691611044
transform 1 0 728 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1691611044
transform 1 0 1972 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_2
timestamp 1691611044
transform 1 0 9166 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_0
timestamp 1691611044
transform 1 0 620 0 1 -672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_1
timestamp 1691611044
transform 1 0 1840 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_2
timestamp 1691611044
transform 1 0 3290 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_3
timestamp 1691611044
transform 1 0 4600 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_4
timestamp 1691611044
transform 1 0 6118 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_5
timestamp 1691611044
transform 1 0 7428 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_6
timestamp 1691611044
transform 1 0 8982 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_7
timestamp 1691611044
transform 1 0 3360 0 1 -1342
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_8
timestamp 1691611044
transform 1 0 4688 0 1 -1342
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_9
timestamp 1691611044
transform 1 0 6218 0 1 -1342
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_10
timestamp 1691611044
transform 1 0 7518 0 1 -1342
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1691611044
transform 1 0 2448 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1691611044
transform 1 0 5278 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1691611044
transform 1 0 8100 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1691611044
transform 1 0 2448 0 1 -670
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1691611044
transform 1 0 2448 0 1 -1342
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1691611044
transform 1 0 5278 0 1 -668
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1691611044
transform 1 0 5278 0 1 -1342
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1691611044
transform 1 0 8100 0 1 -668
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1691611044
transform 1 0 8100 0 1 -1342
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0
timestamp 1691611044
transform 1 0 480 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1691611044
transform 1 0 1714 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_2
timestamp 1691611044
transform 1 0 3228 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_3
timestamp 1691611044
transform 1 0 4528 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_4
timestamp 1691611044
transform 1 0 6038 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_5
timestamp 1691611044
transform 1 0 7348 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_6
timestamp 1691611044
transform 1 0 8890 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_7
timestamp 1691611044
transform 1 0 0 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_8
timestamp 1691611044
transform 1 0 1214 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_9
timestamp 1691611044
transform 1 0 2658 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_10
timestamp 1691611044
transform 1 0 3968 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_11
timestamp 1691611044
transform 1 0 5478 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_12
timestamp 1691611044
transform 1 0 6788 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_13
timestamp 1691611044
transform 1 0 8308 0 1 -1342
box -38 -48 682 592
<< end >>
