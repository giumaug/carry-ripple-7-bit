magic
tech sky130A
magscale 1 2
timestamp 1742633757
<< nwell >>
rect -40 260 9580 592
rect 2540 -100 2710 -78
rect 2540 -400 2630 -100
rect 2540 -420 2710 -400
rect 3234 -409 3270 -88
rect 3870 -409 3937 -88
rect 4543 -409 4568 -88
rect 5185 -406 5245 -88
rect 5394 -398 5460 -86
rect 5394 -406 5580 -398
rect 5185 -407 5580 -406
rect 6045 -407 6090 -86
rect 6700 -407 6754 -86
rect 7365 -407 7395 -86
rect 8013 -407 8068 -86
rect 8200 -90 8370 -80
rect 8200 -400 8300 -90
rect 5188 -410 5580 -407
rect 8200 -410 8370 -400
rect 8895 -407 8952 -86
rect 5400 -760 5570 -750
rect 671 -1081 692 -760
rect 1120 -1081 1182 -760
rect 1880 -1081 1940 -760
rect 2360 -1081 2417 -760
rect 2570 -1080 2630 -760
rect 5400 -1080 5450 -760
rect 2570 -1090 2750 -1080
rect 5400 -1090 5570 -1080
rect 6155 -1081 6184 -760
rect 7460 -1081 7484 -760
rect 8224 -1081 8276 -760
rect 8986 -1081 9131 -760
<< pwell >>
rect 1109 -49 1235 60
rect 1665 -48 1720 48
<< locali >>
rect 454 527 502 561
rect 1121 527 1217 561
rect 1665 527 1719 561
rect 2349 527 2453 561
rect 2532 527 2668 561
rect 3115 527 3233 561
rect 3866 527 3973 561
rect 4427 527 4530 561
rect 5170 527 5282 561
rect 5363 527 5481 561
rect 5928 527 6044 561
rect 6675 527 6792 561
rect 7246 527 7352 561
rect 7990 527 8104 561
rect 8184 527 8313 561
rect 8759 527 8894 561
rect 10 280 90 300
rect 10 240 30 280
rect 70 240 90 280
rect 10 220 90 240
rect 2026 249 2101 260
rect 2026 243 2051 249
rect 2085 243 2101 249
rect 437 -17 504 17
rect 1117 -17 1221 17
rect 1656 -18 1720 17
rect 2348 -17 2457 17
rect 2526 -17 2661 17
rect 3115 -17 3235 17
rect 3863 -17 3973 17
rect 4417 -17 4534 17
rect 5170 -17 5285 17
rect 5359 -17 5483 17
rect 5925 -17 6047 17
rect 6678 -17 6794 17
rect 7237 -17 7354 17
rect 7981 -17 8104 17
rect 8178 -17 8315 17
rect 8768 -17 8894 17
rect 5110 -109 5280 -104
rect 529 -145 624 -111
rect 1169 -145 1231 -109
rect 1756 -143 1842 -109
rect 2388 -143 2452 -109
rect 2523 -143 2664 -109
rect 3208 -143 3316 -109
rect 3828 -143 3974 -109
rect 4513 -143 4604 -109
rect 5110 -120 5282 -109
rect 5149 -141 5282 -120
rect 5367 -141 5487 -107
rect 6027 -141 6121 -107
rect 6655 -141 6799 -107
rect 7337 -141 7433 -107
rect 7977 -141 8103 -107
rect 8183 -141 8314 -107
rect 8857 -141 8987 -107
rect 545 -689 624 -655
rect 1155 -660 1220 -650
rect 5126 -653 5281 -651
rect 1163 -687 1217 -660
rect 1762 -687 1843 -653
rect 2383 -687 2453 -653
rect 2533 -687 2665 -653
rect 3200 -687 3293 -653
rect 3830 -687 3976 -653
rect 4502 -687 4603 -653
rect 5126 -686 5285 -653
rect 5362 -685 5484 -651
rect 6027 -686 6126 -651
rect 6661 -685 6793 -651
rect 7333 -685 7433 -651
rect 7974 -685 8107 -651
rect 8189 -685 8313 -651
rect 8859 -685 8997 -651
rect 5126 -687 5281 -686
rect 626 -815 732 -781
rect 1092 -815 1222 -781
rect 1844 -815 1977 -781
rect 2332 -815 2451 -781
rect 2537 -815 2660 -781
rect 3293 -815 3364 -781
rect 3895 -815 3973 -781
rect 4600 -815 4692 -781
rect 5233 -815 5283 -781
rect 5369 -815 5490 -781
rect 6111 -815 6226 -781
rect 6763 -815 6792 -781
rect 7425 -815 7523 -781
rect 8060 -815 8106 -781
rect 8187 -815 8318 -781
rect 8944 -815 9174 -781
rect 632 -1359 732 -1325
rect 1087 -1359 1224 -1325
rect 1851 -1359 1975 -1325
rect 2330 -1359 2455 -1325
rect 2528 -1359 2666 -1325
rect 3293 -1359 3363 -1325
rect 3902 -1360 3974 -1325
rect 4603 -1359 4694 -1325
rect 5228 -1359 5285 -1325
rect 5368 -1359 5484 -1325
rect 6113 -1359 6225 -1325
rect 6758 -1359 6811 -1325
rect 7426 -1359 7524 -1325
rect 8062 -1359 8110 -1325
rect 8186 -1359 8313 -1325
rect 8945 -1359 9174 -1325
<< viali >>
rect 8680 390 8720 430
rect 30 240 70 280
rect 571 270 606 306
rect 1061 289 1095 323
rect 2295 289 2329 323
rect 3810 290 3850 330
rect 5095 307 5129 341
rect 6600 300 6640 340
rect 210 220 250 260
rect 680 218 716 253
rect 1240 230 1280 270
rect 5880 260 5914 295
rect 7920 290 7960 330
rect 9460 290 9500 330
rect 1429 215 1463 249
rect 1915 215 1950 251
rect 2051 215 2085 249
rect 2690 220 2730 260
rect 2873 223 2907 258
rect 3057 221 3092 255
rect 3320 215 3356 250
rect 3430 210 3470 250
rect 3990 220 4030 260
rect 4181 221 4215 255
rect 4370 200 4404 234
rect 4720 210 4760 250
rect 4865 218 4899 253
rect 5507 223 5541 258
rect 5690 220 5730 260
rect 6240 215 6274 249
rect 6375 215 6409 249
rect 6803 225 6840 260
rect 7001 221 7035 255
rect 7185 209 7219 245
rect 7433 215 7467 249
rect 7550 217 7584 252
rect 8339 221 8373 255
rect 8525 215 8559 249
rect 9092 215 9126 249
rect 9220 210 9260 250
rect 397 153 431 187
rect 1610 140 1650 180
rect 37 -256 71 -220
rect 3994 -260 4034 -220
rect 8334 -290 8370 -251
rect 213 -457 258 -417
rect 480 -457 514 -423
rect 1438 -455 1472 -421
rect 1565 -455 1600 -421
rect 1694 -455 1728 -421
rect 2882 -453 2916 -419
rect 3138 -455 3172 -421
rect 4192 -455 4226 -421
rect 4448 -455 4482 -421
rect 5690 -450 5730 -408
rect 5820 -460 5860 -420
rect 5958 -453 5992 -419
rect 7020 -450 7060 -410
rect 7140 -450 7180 -410
rect 7268 -453 7302 -419
rect 8540 -450 8580 -410
rect 8790 -453 8824 -419
rect 390 -570 430 -530
rect 1251 -575 1285 -541
rect 2680 -560 2720 -520
rect 3055 -580 3090 -543
rect 4360 -570 4400 -530
rect 6810 -570 6850 -530
rect 8706 -567 8741 -533
rect 570 -970 610 -930
rect 1781 -967 1815 -933
rect 3239 -1053 3273 -1019
rect 4540 -1060 4580 -1020
rect 6050 -1050 6090 -1010
rect 8400 -1070 8435 -1036
rect 8890 -1050 8930 -1010
rect 85 -1127 119 -1093
rect 202 -1127 242 -1087
rect 1300 -1140 1340 -1090
rect 1416 -1127 1450 -1093
rect 2747 -1130 2783 -1093
rect 2860 -1127 2894 -1093
rect 4053 -1127 4087 -1093
rect 4170 -1127 4204 -1093
rect 5563 -1127 5597 -1093
rect 5680 -1127 5714 -1093
rect 6873 -1127 6907 -1093
rect 6990 -1127 7024 -1093
rect 8510 -1127 8544 -1093
rect 7289 -1230 7323 -1193
<< metal1 >>
rect 444 496 498 592
rect 1115 496 1218 592
rect 1669 496 1720 592
rect 2354 496 2456 592
rect 2537 496 2661 592
rect 3110 496 3238 592
rect 3851 496 3977 592
rect 4423 496 4532 592
rect 5167 496 5282 592
rect 5367 496 5484 592
rect 5934 496 6044 592
rect 6679 496 6791 592
rect 7240 496 7354 592
rect 7987 496 8105 592
rect 8188 496 8312 592
rect 8765 496 8898 592
rect 8650 450 8740 460
rect 8650 380 8660 450
rect 8730 380 8740 450
rect 8650 370 8740 380
rect 5070 350 5150 360
rect 2270 340 2350 350
rect 1040 330 1120 340
rect 550 306 619 330
rect 10 290 90 300
rect 10 230 20 290
rect 80 230 90 290
rect 10 220 90 230
rect 190 260 270 290
rect 550 270 571 306
rect 606 270 619 306
rect 660 280 740 290
rect 660 270 670 280
rect 550 260 619 270
rect 190 220 210 260
rect 250 220 270 260
rect 190 210 270 220
rect 650 220 670 270
rect 730 270 740 280
rect 1040 270 1050 330
rect 1110 270 1120 330
rect 730 220 760 270
rect 1040 260 1120 270
rect 1200 280 1310 290
rect 2270 280 2280 340
rect 2340 280 2350 340
rect 3780 340 3860 350
rect 3780 280 3790 340
rect 3850 280 3860 340
rect 5070 290 5080 350
rect 5140 290 5150 350
rect 6580 350 6660 360
rect 5860 310 5940 320
rect 5070 280 5150 290
rect 5490 280 5570 290
rect 650 218 680 220
rect 716 218 760 220
rect 650 210 760 218
rect 1200 220 1210 280
rect 1270 270 1310 280
rect 1900 270 1980 280
rect 2270 270 2350 280
rect 2680 270 2760 280
rect 1280 230 1310 270
rect 1270 220 1310 230
rect 1200 210 1310 220
rect 1413 249 1490 270
rect 1413 215 1429 249
rect 1463 215 1490 249
rect 360 190 451 200
rect 1413 190 1490 215
rect 1900 210 1910 270
rect 1970 210 1980 270
rect 2026 250 2100 258
rect 1900 200 1980 210
rect 2020 249 2100 250
rect 2020 240 2051 249
rect 2085 240 2100 249
rect 1590 190 1670 200
rect 360 130 380 190
rect 440 130 451 190
rect 360 120 451 130
rect 1590 130 1600 190
rect 1660 130 1670 190
rect 2020 180 2030 240
rect 2090 180 2100 240
rect 2680 210 2690 270
rect 2750 210 2760 270
rect 2680 200 2760 210
rect 2850 270 2930 280
rect 3410 270 3490 280
rect 3780 270 3860 280
rect 3960 270 4040 280
rect 2850 210 2860 270
rect 2920 210 2930 270
rect 2850 190 2930 210
rect 3050 260 3130 270
rect 3313 260 3362 270
rect 3050 255 3060 260
rect 3050 221 3057 255
rect 3050 200 3060 221
rect 3120 200 3130 260
rect 3050 190 3130 200
rect 3280 250 3362 260
rect 3280 215 3320 250
rect 3356 215 3362 250
rect 3280 199 3362 215
rect 3410 210 3420 270
rect 3480 210 3490 270
rect 3410 200 3490 210
rect 3960 210 3970 270
rect 4030 210 4040 270
rect 4167 260 4235 265
rect 3960 200 4040 210
rect 4160 255 4240 260
rect 4160 250 4181 255
rect 4215 250 4240 255
rect 3280 190 3360 199
rect 4160 190 4170 250
rect 4230 190 4240 250
rect 4160 180 4240 190
rect 4360 250 4440 260
rect 4360 190 4370 250
rect 4430 190 4440 250
rect 4700 210 4720 270
rect 4780 210 4800 270
rect 4700 200 4800 210
rect 4840 260 4920 271
rect 4360 180 4440 190
rect 4840 199 4850 260
rect 4910 199 4920 260
rect 5490 220 5500 280
rect 5560 220 5570 280
rect 5490 210 5570 220
rect 5670 270 5760 280
rect 5670 210 5680 270
rect 5740 210 5760 270
rect 5860 250 5870 310
rect 5930 250 5940 310
rect 6580 290 6590 350
rect 6650 290 6660 350
rect 9440 340 9520 350
rect 6580 280 6660 290
rect 7900 330 7980 340
rect 7520 270 7600 280
rect 6780 260 6860 270
rect 5860 240 5940 250
rect 6200 250 6330 260
rect 2020 170 2100 180
rect 4840 179 4920 199
rect 5670 170 5760 210
rect 6200 190 6220 250
rect 6280 190 6330 250
rect 6200 170 6330 190
rect 6360 250 6440 260
rect 6360 190 6370 250
rect 6430 190 6440 250
rect 6780 200 6790 260
rect 6850 200 6860 260
rect 6780 190 6860 200
rect 6980 260 7060 270
rect 7520 260 7530 270
rect 6980 200 6990 260
rect 7050 200 7060 260
rect 6980 190 7060 200
rect 7170 250 7250 260
rect 7170 190 7180 250
rect 7240 190 7250 250
rect 6360 180 6440 190
rect 7170 180 7250 190
rect 7399 250 7480 260
rect 7399 190 7410 250
rect 7470 190 7480 250
rect 7510 210 7530 260
rect 7590 260 7600 270
rect 7900 270 7910 330
rect 7970 270 7980 330
rect 7900 260 7980 270
rect 8290 290 8380 310
rect 7590 210 7630 260
rect 8290 230 8300 290
rect 8360 270 8380 290
rect 9440 280 9450 340
rect 9510 280 9520 340
rect 8360 255 8399 270
rect 8290 221 8339 230
rect 8373 221 8399 255
rect 8290 210 8399 221
rect 8500 260 8590 270
rect 7520 200 7600 210
rect 8500 200 8510 260
rect 8570 200 8590 260
rect 8500 190 8590 200
rect 9050 260 9180 270
rect 9050 200 9060 260
rect 9120 249 9180 260
rect 9126 215 9180 249
rect 9120 200 9180 215
rect 9050 190 9180 200
rect 9210 260 9310 280
rect 9440 270 9520 280
rect 9210 200 9220 260
rect 9280 200 9310 260
rect 9210 190 9310 200
rect 7399 170 7480 190
rect 1590 120 1670 130
rect 447 -49 518 48
rect 1114 -49 1223 48
rect 1665 -48 1720 48
rect 2352 17 2461 48
rect 2348 -17 2461 17
rect 2352 -49 2461 -17
rect 2535 -48 2666 48
rect 3111 -48 3238 48
rect 3867 -48 3973 48
rect 4423 -14 4532 48
rect 4422 -48 4651 -14
rect 5166 -48 5285 48
rect 5365 -48 5486 48
rect 5933 -48 6045 48
rect 6675 -48 6794 48
rect 7244 -48 7357 48
rect 7986 -48 8108 48
rect 8185 -48 8314 48
rect 8761 -48 8894 48
rect 541 -176 635 -80
rect 1154 -174 1219 -80
rect 1762 -174 1846 -78
rect 2381 -174 2454 -78
rect 2532 -174 2664 -78
rect 3200 -174 3300 -78
rect 3835 -174 3976 -78
rect 4504 -174 4606 -78
rect 5144 -172 5283 -78
rect 5361 -172 5487 -76
rect 6023 -172 6124 -76
rect 6665 -172 6794 -76
rect 7334 -172 7431 -76
rect 7974 -172 8104 -76
rect 8186 -172 8313 -76
rect 8845 -172 8988 -76
rect 20 -220 100 -210
rect 20 -280 30 -220
rect 90 -280 100 -220
rect 20 -290 100 -280
rect 3980 -220 4060 -210
rect 3980 -280 3990 -220
rect 4050 -280 4060 -220
rect 3980 -290 4060 -280
rect 8310 -230 8390 -220
rect 8310 -290 8320 -230
rect 8380 -290 8390 -230
rect 8310 -300 8390 -290
rect 180 -400 260 -390
rect 180 -460 190 -400
rect 250 -417 270 -400
rect 258 -457 270 -417
rect 250 -460 270 -457
rect 180 -470 270 -460
rect 470 -423 550 -390
rect 1420 -400 1500 -390
rect 1420 -405 1430 -400
rect 470 -457 480 -423
rect 514 -457 550 -423
rect 470 -470 550 -457
rect 1417 -460 1430 -405
rect 1490 -405 1500 -400
rect 1550 -400 1630 -380
rect 2850 -390 2930 -380
rect 1490 -460 1509 -405
rect 1417 -468 1509 -460
rect 1550 -460 1560 -400
rect 1620 -460 1630 -400
rect 1420 -470 1500 -468
rect 1550 -470 1630 -460
rect 1680 -400 1760 -390
rect 1680 -460 1690 -400
rect 1750 -460 1760 -400
rect 2850 -450 2860 -390
rect 2920 -450 2930 -390
rect 2850 -453 2882 -450
rect 2916 -453 2930 -450
rect 2850 -460 2930 -453
rect 3130 -400 3210 -390
rect 3130 -421 3140 -400
rect 3130 -455 3138 -421
rect 3130 -460 3140 -455
rect 3200 -460 3210 -400
rect 1680 -470 1760 -460
rect 3130 -470 3210 -460
rect 4170 -400 4250 -390
rect 4170 -460 4180 -400
rect 4240 -460 4250 -400
rect 4170 -470 4250 -460
rect 4440 -400 4520 -390
rect 4440 -421 4450 -400
rect 4440 -455 4448 -421
rect 4440 -460 4450 -455
rect 4510 -460 4520 -400
rect 5670 -408 5750 -380
rect 5670 -450 5690 -408
rect 5730 -450 5750 -408
rect 5670 -460 5750 -450
rect 5800 -400 5880 -390
rect 5800 -460 5810 -400
rect 5870 -460 5880 -400
rect 4440 -470 4520 -460
rect 5800 -470 5880 -460
rect 5940 -399 6020 -390
rect 5940 -460 5950 -399
rect 6010 -460 6020 -399
rect 5940 -470 6020 -460
rect 6990 -400 7070 -390
rect 6990 -460 7000 -400
rect 7060 -460 7070 -400
rect 6990 -470 7070 -460
rect 7120 -400 7200 -390
rect 7120 -460 7130 -400
rect 7190 -460 7200 -400
rect 7120 -470 7200 -460
rect 7260 -400 7340 -390
rect 7260 -419 7270 -400
rect 7260 -453 7268 -419
rect 7260 -460 7270 -453
rect 7330 -460 7340 -400
rect 7260 -470 7340 -460
rect 8520 -400 8600 -390
rect 8520 -460 8530 -400
rect 8590 -460 8600 -400
rect 8520 -470 8600 -460
rect 8780 -410 8860 -400
rect 8780 -470 8790 -410
rect 8850 -470 8860 -410
rect 8780 -480 8860 -470
rect 2650 -510 2730 -500
rect 8670 -510 8750 -500
rect 380 -520 460 -510
rect 380 -580 390 -520
rect 450 -580 460 -520
rect 380 -590 460 -580
rect 1220 -520 1300 -510
rect 1220 -580 1230 -520
rect 1290 -580 1300 -520
rect 2650 -570 2660 -510
rect 2720 -570 2730 -510
rect 2650 -580 2730 -570
rect 3030 -520 3110 -510
rect 3030 -580 3040 -520
rect 3100 -580 3110 -520
rect 1220 -590 1300 -580
rect 3030 -590 3110 -580
rect 4330 -520 4410 -510
rect 4330 -580 4340 -520
rect 4400 -580 4410 -520
rect 4330 -590 4410 -580
rect 6780 -520 6860 -510
rect 6780 -580 6790 -520
rect 6850 -580 6860 -520
rect 8670 -570 8680 -510
rect 8740 -533 8750 -510
rect 8741 -567 8750 -533
rect 8740 -570 8750 -567
rect 8670 -580 8750 -570
rect 6780 -590 6860 -580
rect 537 -720 623 -624
rect 1167 -718 1217 -624
rect 1755 -718 1843 -622
rect 2386 -718 2453 -622
rect 2535 -718 2666 -622
rect 3204 -718 3295 -622
rect 3834 -718 3976 -622
rect 4515 -718 4604 -622
rect 5144 -720 5283 -620
rect 5365 -716 5487 -620
rect 6024 -716 6125 -620
rect 6666 -716 6795 -620
rect 7336 -716 7436 -620
rect 7977 -716 8107 -620
rect 8186 -716 8315 -620
rect 8856 -716 8992 -620
rect 634 -846 735 -750
rect 1086 -846 1219 -750
rect 1851 -846 1983 -750
rect 2335 -846 2454 -750
rect 2535 -846 2662 -750
rect 3298 -846 3364 -750
rect 3902 -846 3974 -750
rect 4606 -846 4693 -750
rect 5232 -846 5284 -750
rect 5366 -846 5484 -750
rect 6116 -846 6225 -750
rect 6756 -846 6806 -750
rect 7424 -846 7523 -750
rect 8065 -846 8112 -750
rect 8181 -846 8314 -750
rect 8937 -846 9175 -750
rect 560 -920 640 -910
rect 560 -980 570 -920
rect 630 -980 640 -920
rect 560 -990 640 -980
rect 1770 -920 1850 -910
rect 1770 -980 1779 -920
rect 1839 -980 1850 -920
rect 1770 -990 1850 -980
rect 6030 -970 6050 -910
rect 6110 -970 6120 -910
rect 3220 -1000 3300 -990
rect 3220 -1060 3230 -1000
rect 3290 -1060 3300 -1000
rect 4520 -1000 4600 -990
rect 4520 -1060 4530 -1000
rect 4590 -1060 4600 -1000
rect 6030 -1010 6120 -970
rect 8870 -1000 8950 -990
rect 6030 -1050 6050 -1010
rect 6090 -1050 6120 -1010
rect 180 -1070 260 -1060
rect 2840 -1070 2920 -1060
rect 3220 -1070 3300 -1060
rect 4020 -1070 4100 -1060
rect 59 -1080 140 -1070
rect 59 -1140 70 -1080
rect 130 -1140 140 -1080
rect 180 -1130 190 -1070
rect 250 -1130 260 -1070
rect 1400 -1080 1480 -1070
rect 180 -1140 260 -1130
rect 1280 -1090 1360 -1080
rect 1280 -1140 1300 -1090
rect 1340 -1140 1360 -1090
rect 59 -1150 140 -1140
rect 1280 -1160 1360 -1140
rect 1400 -1140 1410 -1080
rect 1470 -1140 1480 -1080
rect 1400 -1150 1480 -1140
rect 2720 -1080 2800 -1070
rect 2720 -1140 2730 -1080
rect 2790 -1140 2800 -1080
rect 2840 -1130 2850 -1070
rect 2910 -1130 2920 -1070
rect 2840 -1140 2920 -1130
rect 4020 -1130 4030 -1070
rect 4090 -1130 4100 -1070
rect 4020 -1140 4100 -1130
rect 4150 -1070 4230 -1060
rect 4520 -1070 4600 -1060
rect 5670 -1070 5750 -1060
rect 6030 -1070 6120 -1050
rect 8370 -1010 8450 -1000
rect 8370 -1070 8380 -1010
rect 8440 -1070 8450 -1010
rect 8870 -1060 8880 -1000
rect 8940 -1060 8950 -1000
rect 4150 -1130 4160 -1070
rect 4220 -1130 4230 -1070
rect 4150 -1140 4230 -1130
rect 5540 -1080 5620 -1070
rect 5540 -1140 5550 -1080
rect 5610 -1140 5620 -1080
rect 5670 -1130 5680 -1070
rect 5740 -1130 5750 -1070
rect 5670 -1140 5750 -1130
rect 6850 -1080 6930 -1070
rect 6850 -1140 6860 -1080
rect 6920 -1140 6930 -1080
rect 2720 -1150 2800 -1140
rect 5540 -1150 5620 -1140
rect 6850 -1150 6930 -1140
rect 6970 -1080 7050 -1070
rect 8370 -1080 8450 -1070
rect 8490 -1070 8570 -1060
rect 8870 -1070 8950 -1060
rect 6970 -1140 6980 -1080
rect 7040 -1140 7050 -1080
rect 8490 -1130 8500 -1070
rect 8560 -1130 8570 -1070
rect 8490 -1140 8570 -1130
rect 6970 -1150 7050 -1140
rect 7270 -1170 7360 -1160
rect 7270 -1193 7290 -1170
rect 7270 -1230 7289 -1193
rect 7350 -1230 7360 -1170
rect 7270 -1240 7360 -1230
rect 7270 -1250 7309 -1240
rect 637 -1390 734 -1294
rect 1090 -1390 1222 -1294
rect 1854 -1390 1980 -1294
rect 2336 -1390 2454 -1294
rect 2534 -1390 2665 -1294
rect 3297 -1390 3364 -1294
rect 3906 -1390 3978 -1294
rect 4606 -1390 4696 -1294
rect 5233 -1390 5292 -1294
rect 5364 -1390 5488 -1294
rect 6116 -1390 6226 -1294
rect 6765 -1390 6813 -1294
rect 7425 -1390 7527 -1294
rect 8065 -1390 8105 -1294
rect 8188 -1390 8316 -1294
rect 8944 -1390 9170 -1294
<< via1 >>
rect 8660 430 8730 450
rect 8660 390 8680 430
rect 8680 390 8720 430
rect 8720 390 8730 430
rect 8660 380 8730 390
rect 20 280 80 290
rect 20 240 30 280
rect 30 240 70 280
rect 70 240 80 280
rect 20 230 80 240
rect 670 253 730 280
rect 1050 323 1110 330
rect 1050 289 1061 323
rect 1061 289 1095 323
rect 1095 289 1110 323
rect 1050 270 1110 289
rect 670 220 680 253
rect 680 220 716 253
rect 716 220 730 253
rect 2280 323 2340 340
rect 2280 289 2295 323
rect 2295 289 2329 323
rect 2329 289 2340 323
rect 2280 280 2340 289
rect 3790 330 3850 340
rect 3790 290 3810 330
rect 3810 290 3850 330
rect 3790 280 3850 290
rect 5080 341 5140 350
rect 5080 307 5095 341
rect 5095 307 5129 341
rect 5129 307 5140 341
rect 5080 290 5140 307
rect 1210 270 1270 280
rect 1210 230 1240 270
rect 1240 230 1270 270
rect 1210 220 1270 230
rect 1910 251 1970 270
rect 1910 215 1915 251
rect 1915 215 1950 251
rect 1950 215 1970 251
rect 1910 210 1970 215
rect 380 187 440 190
rect 380 153 397 187
rect 397 153 431 187
rect 431 153 440 187
rect 380 130 440 153
rect 1600 180 1660 190
rect 1600 140 1610 180
rect 1610 140 1650 180
rect 1650 140 1660 180
rect 1600 130 1660 140
rect 2030 215 2051 240
rect 2051 215 2085 240
rect 2085 215 2090 240
rect 2030 180 2090 215
rect 2690 260 2750 270
rect 2690 220 2730 260
rect 2730 220 2750 260
rect 2690 210 2750 220
rect 2860 258 2920 270
rect 2860 223 2873 258
rect 2873 223 2907 258
rect 2907 223 2920 258
rect 2860 210 2920 223
rect 3060 255 3120 260
rect 3060 221 3092 255
rect 3092 221 3120 255
rect 3060 200 3120 221
rect 3420 250 3480 270
rect 3420 210 3430 250
rect 3430 210 3470 250
rect 3470 210 3480 250
rect 3970 260 4030 270
rect 3970 220 3990 260
rect 3990 220 4030 260
rect 3970 210 4030 220
rect 4170 221 4181 250
rect 4181 221 4215 250
rect 4215 221 4230 250
rect 4170 190 4230 221
rect 4370 234 4430 250
rect 4370 200 4404 234
rect 4404 200 4430 234
rect 4370 190 4430 200
rect 4720 250 4780 270
rect 4720 210 4760 250
rect 4760 210 4780 250
rect 4850 253 4910 260
rect 4850 218 4865 253
rect 4865 218 4899 253
rect 4899 218 4910 253
rect 4850 199 4910 218
rect 5500 258 5560 280
rect 5500 223 5507 258
rect 5507 223 5541 258
rect 5541 223 5560 258
rect 5500 220 5560 223
rect 5680 260 5740 270
rect 5680 220 5690 260
rect 5690 220 5730 260
rect 5730 220 5740 260
rect 5680 210 5740 220
rect 5870 295 5930 310
rect 5870 260 5880 295
rect 5880 260 5914 295
rect 5914 260 5930 295
rect 5870 250 5930 260
rect 6590 340 6650 350
rect 6590 300 6600 340
rect 6600 300 6640 340
rect 6640 300 6650 340
rect 6590 290 6650 300
rect 6220 249 6280 250
rect 6220 215 6240 249
rect 6240 215 6274 249
rect 6274 215 6280 249
rect 6220 190 6280 215
rect 6370 249 6430 250
rect 6370 215 6375 249
rect 6375 215 6409 249
rect 6409 215 6430 249
rect 6370 190 6430 215
rect 6790 225 6803 260
rect 6803 225 6840 260
rect 6840 225 6850 260
rect 6790 200 6850 225
rect 6990 255 7050 260
rect 6990 221 7001 255
rect 7001 221 7035 255
rect 7035 221 7050 255
rect 6990 200 7050 221
rect 7180 245 7240 250
rect 7180 209 7185 245
rect 7185 209 7219 245
rect 7219 209 7240 245
rect 7180 190 7240 209
rect 7410 249 7470 250
rect 7410 215 7433 249
rect 7433 215 7467 249
rect 7467 215 7470 249
rect 7410 190 7470 215
rect 7530 252 7590 270
rect 7910 290 7920 330
rect 7920 290 7960 330
rect 7960 290 7970 330
rect 7910 270 7970 290
rect 7530 217 7550 252
rect 7550 217 7584 252
rect 7584 217 7590 252
rect 7530 210 7590 217
rect 8300 255 8360 290
rect 9450 330 9510 340
rect 9450 290 9460 330
rect 9460 290 9500 330
rect 9500 290 9510 330
rect 9450 280 9510 290
rect 8300 230 8339 255
rect 8339 230 8360 255
rect 8510 249 8570 260
rect 8510 215 8525 249
rect 8525 215 8559 249
rect 8559 215 8570 249
rect 8510 200 8570 215
rect 9060 249 9120 260
rect 9060 215 9092 249
rect 9092 215 9120 249
rect 9060 200 9120 215
rect 9220 250 9280 260
rect 9220 210 9260 250
rect 9260 210 9280 250
rect 9220 200 9280 210
rect 30 -256 37 -220
rect 37 -256 71 -220
rect 71 -256 90 -220
rect 30 -280 90 -256
rect 3990 -260 3994 -220
rect 3994 -260 4034 -220
rect 4034 -260 4050 -220
rect 3990 -280 4050 -260
rect 8320 -251 8380 -230
rect 8320 -290 8334 -251
rect 8334 -290 8370 -251
rect 8370 -290 8380 -251
rect 190 -417 250 -400
rect 190 -457 213 -417
rect 213 -457 250 -417
rect 190 -460 250 -457
rect 1430 -421 1490 -400
rect 1430 -455 1438 -421
rect 1438 -455 1472 -421
rect 1472 -455 1490 -421
rect 1430 -460 1490 -455
rect 1560 -421 1620 -400
rect 1560 -455 1565 -421
rect 1565 -455 1600 -421
rect 1600 -455 1620 -421
rect 1560 -460 1620 -455
rect 1690 -421 1750 -400
rect 1690 -455 1694 -421
rect 1694 -455 1728 -421
rect 1728 -455 1750 -421
rect 1690 -460 1750 -455
rect 2860 -419 2920 -390
rect 2860 -450 2882 -419
rect 2882 -450 2916 -419
rect 2916 -450 2920 -419
rect 3140 -421 3200 -400
rect 3140 -455 3172 -421
rect 3172 -455 3200 -421
rect 3140 -460 3200 -455
rect 4180 -421 4240 -400
rect 4180 -455 4192 -421
rect 4192 -455 4226 -421
rect 4226 -455 4240 -421
rect 4180 -460 4240 -455
rect 4450 -421 4510 -400
rect 4450 -455 4482 -421
rect 4482 -455 4510 -421
rect 4450 -460 4510 -455
rect 5810 -420 5870 -400
rect 5810 -460 5820 -420
rect 5820 -460 5860 -420
rect 5860 -460 5870 -420
rect 5950 -419 6010 -399
rect 5950 -453 5958 -419
rect 5958 -453 5992 -419
rect 5992 -453 6010 -419
rect 5950 -460 6010 -453
rect 7000 -410 7060 -400
rect 7000 -450 7020 -410
rect 7020 -450 7060 -410
rect 7000 -460 7060 -450
rect 7130 -410 7190 -400
rect 7130 -450 7140 -410
rect 7140 -450 7180 -410
rect 7180 -450 7190 -410
rect 7130 -460 7190 -450
rect 7270 -419 7330 -400
rect 7270 -453 7302 -419
rect 7302 -453 7330 -419
rect 7270 -460 7330 -453
rect 8530 -410 8590 -400
rect 8530 -450 8540 -410
rect 8540 -450 8580 -410
rect 8580 -450 8590 -410
rect 8530 -460 8590 -450
rect 8790 -419 8850 -410
rect 8790 -453 8824 -419
rect 8824 -453 8850 -419
rect 8790 -470 8850 -453
rect 390 -530 450 -520
rect 390 -570 430 -530
rect 430 -570 450 -530
rect 390 -580 450 -570
rect 1230 -541 1290 -520
rect 1230 -575 1251 -541
rect 1251 -575 1285 -541
rect 1285 -575 1290 -541
rect 1230 -580 1290 -575
rect 2660 -520 2720 -510
rect 2660 -560 2680 -520
rect 2680 -560 2720 -520
rect 2660 -570 2720 -560
rect 3040 -543 3100 -520
rect 3040 -580 3055 -543
rect 3055 -580 3090 -543
rect 3090 -580 3100 -543
rect 4340 -530 4400 -520
rect 4340 -570 4360 -530
rect 4360 -570 4400 -530
rect 4340 -580 4400 -570
rect 6790 -530 6850 -520
rect 6790 -570 6810 -530
rect 6810 -570 6850 -530
rect 6790 -580 6850 -570
rect 8680 -533 8740 -510
rect 8680 -567 8706 -533
rect 8706 -567 8740 -533
rect 8680 -570 8740 -567
rect 570 -930 630 -920
rect 570 -970 610 -930
rect 610 -970 630 -930
rect 570 -980 630 -970
rect 1779 -933 1839 -920
rect 1779 -967 1781 -933
rect 1781 -967 1815 -933
rect 1815 -967 1839 -933
rect 1779 -980 1839 -967
rect 6050 -970 6110 -910
rect 3230 -1019 3290 -1000
rect 3230 -1053 3239 -1019
rect 3239 -1053 3273 -1019
rect 3273 -1053 3290 -1019
rect 3230 -1060 3290 -1053
rect 4530 -1020 4590 -1000
rect 4530 -1060 4540 -1020
rect 4540 -1060 4580 -1020
rect 4580 -1060 4590 -1020
rect 70 -1093 130 -1080
rect 70 -1127 85 -1093
rect 85 -1127 119 -1093
rect 119 -1127 130 -1093
rect 70 -1140 130 -1127
rect 190 -1087 250 -1070
rect 190 -1127 202 -1087
rect 202 -1127 242 -1087
rect 242 -1127 250 -1087
rect 190 -1130 250 -1127
rect 1410 -1093 1470 -1080
rect 1410 -1127 1416 -1093
rect 1416 -1127 1450 -1093
rect 1450 -1127 1470 -1093
rect 1410 -1140 1470 -1127
rect 2730 -1093 2790 -1080
rect 2730 -1130 2747 -1093
rect 2747 -1130 2783 -1093
rect 2783 -1130 2790 -1093
rect 2730 -1140 2790 -1130
rect 2850 -1093 2910 -1070
rect 2850 -1127 2860 -1093
rect 2860 -1127 2894 -1093
rect 2894 -1127 2910 -1093
rect 2850 -1130 2910 -1127
rect 4030 -1093 4090 -1070
rect 4030 -1127 4053 -1093
rect 4053 -1127 4087 -1093
rect 4087 -1127 4090 -1093
rect 4030 -1130 4090 -1127
rect 8380 -1036 8440 -1010
rect 8380 -1070 8400 -1036
rect 8400 -1070 8435 -1036
rect 8435 -1070 8440 -1036
rect 8880 -1010 8940 -1000
rect 8880 -1050 8890 -1010
rect 8890 -1050 8930 -1010
rect 8930 -1050 8940 -1010
rect 8880 -1060 8940 -1050
rect 4160 -1093 4220 -1070
rect 4160 -1127 4170 -1093
rect 4170 -1127 4204 -1093
rect 4204 -1127 4220 -1093
rect 4160 -1130 4220 -1127
rect 5550 -1093 5610 -1080
rect 5550 -1127 5563 -1093
rect 5563 -1127 5597 -1093
rect 5597 -1127 5610 -1093
rect 5550 -1140 5610 -1127
rect 5680 -1093 5740 -1070
rect 5680 -1127 5714 -1093
rect 5714 -1127 5740 -1093
rect 5680 -1130 5740 -1127
rect 6860 -1093 6920 -1080
rect 6860 -1127 6873 -1093
rect 6873 -1127 6907 -1093
rect 6907 -1127 6920 -1093
rect 6860 -1140 6920 -1127
rect 6980 -1093 7040 -1080
rect 6980 -1127 6990 -1093
rect 6990 -1127 7024 -1093
rect 7024 -1127 7040 -1093
rect 6980 -1140 7040 -1127
rect 8500 -1093 8560 -1070
rect 8500 -1127 8510 -1093
rect 8510 -1127 8544 -1093
rect 8544 -1127 8560 -1093
rect 8500 -1130 8560 -1127
rect 7290 -1193 7350 -1170
rect 7290 -1230 7323 -1193
rect 7323 -1230 7350 -1193
<< metal2 >>
rect 2680 500 2760 530
rect 0 440 100 460
rect 0 380 20 440
rect 80 380 100 440
rect 0 360 100 380
rect 660 440 740 460
rect 720 380 740 440
rect 10 290 90 360
rect 10 230 20 290
rect 80 230 90 290
rect 10 220 90 230
rect 190 180 270 290
rect 180 160 270 180
rect 180 100 190 160
rect 250 100 270 160
rect 360 190 450 200
rect 360 130 380 190
rect 440 130 450 190
rect 550 180 630 330
rect 660 280 740 380
rect 1190 440 1280 460
rect 1190 380 1210 440
rect 1270 380 1280 440
rect 1190 360 1280 380
rect 660 220 670 280
rect 730 220 740 280
rect 1040 330 1120 340
rect 1040 270 1050 330
rect 1110 270 1120 330
rect 1040 260 1120 270
rect 1200 280 1280 360
rect 1900 430 1990 460
rect 1900 370 1910 430
rect 1970 370 1990 430
rect 1900 290 1990 370
rect 2680 440 2690 500
rect 2750 440 2760 500
rect 660 210 740 220
rect 1200 220 1210 280
rect 1270 220 1280 280
rect 1890 270 1990 290
rect 2270 340 2350 350
rect 2270 280 2280 340
rect 2340 280 2350 340
rect 2270 270 2350 280
rect 2680 270 2760 440
rect 3410 500 3490 530
rect 3410 440 3420 500
rect 3480 440 3490 500
rect 8290 500 8380 510
rect 5490 460 5570 480
rect 1200 210 1280 220
rect 360 120 450 130
rect 540 160 630 180
rect 1413 170 1490 270
rect 1890 210 1910 270
rect 1970 210 1990 270
rect 180 80 270 100
rect 380 20 440 120
rect 540 100 560 160
rect 620 100 630 160
rect 540 80 630 100
rect 1390 150 1490 170
rect 1390 90 1410 150
rect 1470 90 1490 150
rect 1390 70 1490 90
rect 1590 190 1670 200
rect 1890 190 1990 210
rect 2020 240 2100 250
rect 1590 130 1600 190
rect 1660 130 1670 190
rect 180 10 260 20
rect 180 -50 190 10
rect 250 -50 260 10
rect 180 -60 260 -50
rect 360 10 440 20
rect 360 -50 370 10
rect 430 -50 440 10
rect 360 -60 440 -50
rect 1420 -60 1500 -50
rect 20 -220 100 -210
rect 20 -280 30 -220
rect 90 -280 100 -220
rect 20 -290 100 -280
rect 180 -370 240 -60
rect 1420 -120 1430 -60
rect 1490 -120 1500 -60
rect 180 -400 260 -370
rect 180 -460 190 -400
rect 250 -460 260 -400
rect 180 -468 260 -460
rect 470 -400 550 -390
rect 530 -460 550 -400
rect 470 -470 550 -460
rect 1420 -400 1500 -120
rect 1590 -60 1670 130
rect 2020 180 2030 240
rect 2090 180 2100 240
rect 2680 210 2690 270
rect 2750 210 2760 270
rect 2680 200 2760 210
rect 2850 270 2930 279
rect 2850 210 2860 270
rect 2920 210 2930 270
rect 2020 141 2100 180
rect 2080 80 2100 141
rect 2020 69 2100 80
rect 2850 100 2930 210
rect 3040 270 3140 280
rect 3040 190 3050 270
rect 3130 190 3140 270
rect 3410 270 3490 440
rect 3960 430 4040 450
rect 3960 370 3970 430
rect 4030 370 4040 430
rect 3780 340 3860 350
rect 3780 280 3790 340
rect 3850 280 3860 340
rect 3780 270 3860 280
rect 3960 270 4040 370
rect 4720 420 4800 430
rect 4720 360 4730 420
rect 4790 360 4800 420
rect 5490 400 5510 460
rect 4720 270 4800 360
rect 5070 350 5150 360
rect 5070 290 5080 350
rect 5140 290 5150 350
rect 5070 280 5150 290
rect 5490 280 5570 400
rect 6150 450 6300 480
rect 6150 390 6220 450
rect 6280 390 6300 450
rect 6150 370 6300 390
rect 5860 310 5940 320
rect 3040 180 3140 190
rect 2850 40 2860 100
rect 2920 40 2930 100
rect 2850 20 2930 40
rect 3280 100 3360 260
rect 3410 210 3420 270
rect 3480 210 3490 270
rect 3410 200 3490 210
rect 3960 210 3970 270
rect 4030 210 4040 270
rect 3960 200 4040 210
rect 4160 250 4240 260
rect 3280 40 3290 100
rect 3350 40 3360 100
rect 3280 20 3360 40
rect 4160 190 4170 250
rect 4230 211 4240 250
rect 4360 250 4440 260
rect 4230 190 4241 211
rect 4160 121 4241 190
rect 4160 60 4170 121
rect 4230 60 4241 121
rect 4160 39 4241 60
rect 4360 190 4370 250
rect 4430 190 4440 250
rect 4700 210 4720 270
rect 4780 210 4800 270
rect 4700 200 4800 210
rect 4839 260 4920 269
rect 1590 -120 1600 -60
rect 1660 -120 1670 -60
rect 1590 -130 1670 -120
rect 4170 -30 4250 -20
rect 4170 -90 4180 -30
rect 4240 -90 4250 -30
rect 1550 -210 1630 -200
rect 1550 -270 1560 -210
rect 1620 -270 1630 -210
rect 3980 -220 4060 -210
rect 1550 -280 1630 -270
rect 2820 -230 2920 -220
rect 1560 -380 1620 -280
rect 2820 -310 2830 -230
rect 2910 -240 2920 -230
rect 2910 -310 2930 -240
rect 3980 -280 3990 -220
rect 4050 -280 4060 -220
rect 3980 -290 4060 -280
rect 2820 -320 2930 -310
rect 1420 -460 1430 -400
rect 1490 -460 1500 -400
rect 1420 -470 1500 -460
rect 1550 -400 1630 -380
rect 2850 -390 2930 -320
rect 1550 -460 1560 -400
rect 1620 -460 1630 -400
rect 1550 -470 1630 -460
rect 1680 -400 1760 -390
rect 1680 -460 1690 -400
rect 1750 -460 1760 -400
rect 2850 -450 2860 -390
rect 2920 -450 2930 -390
rect 2850 -460 2930 -450
rect 3120 -390 3220 -380
rect 1680 -470 1760 -460
rect 3120 -470 3130 -390
rect 3210 -470 3220 -390
rect 4170 -400 4250 -90
rect 4360 -30 4440 190
rect 4839 199 4850 260
rect 4910 199 4920 260
rect 5490 220 5500 280
rect 5560 220 5570 280
rect 5490 210 5570 220
rect 5670 270 5750 280
rect 5670 210 5680 270
rect 5740 210 5750 270
rect 5860 250 5870 310
rect 5930 250 5940 310
rect 6220 260 6300 370
rect 6780 450 6860 470
rect 6780 390 6790 450
rect 6850 390 6860 450
rect 6580 350 6660 360
rect 6580 290 6590 350
rect 6650 290 6660 350
rect 6580 280 6660 290
rect 6780 260 6860 390
rect 7520 440 7600 470
rect 7520 380 7530 440
rect 7590 380 7600 440
rect 7520 270 7600 380
rect 8290 440 8300 500
rect 8360 440 8380 500
rect 9030 500 9130 510
rect 5860 240 5940 250
rect 6190 250 6330 260
rect 4839 140 4920 199
rect 4810 119 4920 140
rect 4810 60 4840 119
rect 4900 60 4920 119
rect 4810 40 4920 60
rect 5670 130 5750 210
rect 6190 190 6220 250
rect 6280 190 6330 250
rect 6190 170 6330 190
rect 6360 250 6440 260
rect 6360 190 6370 250
rect 6430 190 6440 250
rect 6780 200 6790 260
rect 6850 200 6860 260
rect 6780 190 6860 200
rect 6980 260 7059 270
rect 6980 200 6990 260
rect 7050 200 7059 260
rect 6360 130 6440 190
rect 5670 120 5790 130
rect 5670 60 5690 120
rect 5750 60 5790 120
rect 4810 39 4840 40
rect 5670 30 5790 60
rect 6339 100 6440 130
rect 6339 40 6370 100
rect 6430 40 6440 100
rect 6339 30 6440 40
rect 6980 90 7059 200
rect 7170 250 7250 260
rect 7170 190 7180 250
rect 7240 190 7250 250
rect 7170 180 7250 190
rect 7399 250 7480 260
rect 7399 190 7410 250
rect 7470 190 7480 250
rect 7520 210 7530 270
rect 7590 210 7600 270
rect 7900 330 7980 340
rect 7900 270 7910 330
rect 7970 270 7980 330
rect 7900 260 7980 270
rect 8290 290 8380 440
rect 8290 230 8300 290
rect 8360 230 8380 290
rect 8650 450 8740 460
rect 8650 380 8660 450
rect 8730 380 8740 450
rect 9030 420 9040 500
rect 9120 420 9130 500
rect 9030 410 9130 420
rect 8650 370 8740 380
rect 8290 210 8380 230
rect 8500 260 8580 270
rect 7520 200 7600 210
rect 8500 200 8510 260
rect 8570 200 8580 260
rect 7399 170 7480 190
rect 8500 180 8580 200
rect 7400 120 7480 170
rect 8480 130 8580 180
rect 6980 30 6990 90
rect 7050 30 7059 90
rect 6980 20 7059 30
rect 7380 100 7490 120
rect 7380 40 7410 100
rect 7470 40 7490 100
rect 8480 70 8500 130
rect 8560 70 8580 130
rect 8480 50 8580 70
rect 7380 20 7490 40
rect 4360 -90 4370 -30
rect 4430 -90 4440 -30
rect 8310 -40 8390 -30
rect 4360 -100 4440 -90
rect 7120 -80 7200 -70
rect 7120 -140 7130 -80
rect 7190 -140 7200 -80
rect 5800 -220 5880 -210
rect 5800 -280 5810 -220
rect 5870 -280 5880 -220
rect 4170 -460 4180 -400
rect 4240 -460 4250 -400
rect 4170 -470 4250 -460
rect 4440 -400 4520 -390
rect 4440 -460 4450 -400
rect 4510 -460 4520 -400
rect 4440 -470 4520 -460
rect 3120 -480 3220 -470
rect 2650 -510 2730 -498
rect 380 -520 470 -510
rect 380 -580 390 -520
rect 450 -570 470 -520
rect 380 -630 400 -580
rect 460 -630 470 -570
rect 1220 -520 1300 -510
rect 1220 -620 1230 -520
rect 1290 -620 1300 -520
rect 1220 -630 1300 -620
rect 2650 -570 2660 -510
rect 2720 -570 2730 -510
rect 380 -640 470 -630
rect 2650 -710 2730 -570
rect 3030 -520 3110 -510
rect 3030 -620 3040 -520
rect 3100 -620 3110 -520
rect 4330 -520 4410 -510
rect 4330 -580 4340 -520
rect 4400 -580 4410 -520
rect 2650 -770 2660 -710
rect 2720 -770 2730 -710
rect 2650 -780 2730 -770
rect 4330 -710 4410 -580
rect 4330 -770 4340 -710
rect 4400 -770 4410 -710
rect 820 -910 900 -870
rect 2020 -910 2120 -890
rect 560 -920 900 -910
rect 60 -950 140 -940
rect 60 -1010 70 -950
rect 130 -1010 140 -950
rect 560 -980 570 -920
rect 630 -980 900 -920
rect 560 -990 900 -980
rect 1769 -920 2120 -910
rect 1769 -980 1779 -920
rect 1839 -980 2120 -920
rect 1769 -990 2120 -980
rect 2720 -900 2820 -890
rect 2720 -980 2730 -900
rect 2810 -980 2820 -900
rect 2720 -990 2820 -980
rect 60 -1080 140 -1010
rect 60 -1140 70 -1080
rect 130 -1140 140 -1080
rect 60 -1150 140 -1140
rect 180 -1070 260 -1060
rect 180 -1180 190 -1070
rect 250 -1180 260 -1070
rect 1390 -1070 1490 -1060
rect 1280 -1160 1360 -1080
rect 1390 -1150 1400 -1070
rect 1480 -1150 1490 -1070
rect 2720 -1080 2800 -990
rect 3220 -1000 3690 -990
rect 2720 -1140 2730 -1080
rect 2790 -1140 2800 -1080
rect 2720 -1150 2800 -1140
rect 2830 -1060 2930 -1050
rect 2830 -1140 2840 -1060
rect 2920 -1140 2930 -1060
rect 3220 -1060 3230 -1000
rect 3290 -1060 3690 -1000
rect 4330 -1060 4410 -770
rect 5540 -660 5620 -650
rect 5540 -720 5550 -660
rect 5610 -720 5620 -660
rect 3220 -1070 3690 -1060
rect 3610 -1130 3620 -1070
rect 3680 -1130 3690 -1070
rect 3610 -1140 3690 -1130
rect 4020 -1070 4100 -1060
rect 4020 -1130 4030 -1070
rect 4090 -1130 4100 -1070
rect 2830 -1150 2930 -1140
rect 1390 -1160 1490 -1150
rect 180 -1190 260 -1180
rect 1290 -1220 1350 -1160
rect 4020 -1210 4100 -1130
rect 4150 -1070 4410 -1060
rect 4520 -1000 4840 -990
rect 4520 -1060 4530 -1000
rect 4590 -1060 4770 -1000
rect 4830 -1060 4840 -1000
rect 4520 -1070 4840 -1060
rect 4150 -1130 4160 -1070
rect 4220 -1130 4410 -1070
rect 4150 -1140 4410 -1130
rect 5540 -1080 5620 -720
rect 5670 -870 5750 -380
rect 5800 -400 5880 -280
rect 6990 -250 7070 -240
rect 6990 -310 7000 -250
rect 7060 -310 7070 -250
rect 5800 -460 5810 -400
rect 5870 -460 5880 -400
rect 5800 -660 5880 -460
rect 5940 -399 6020 -390
rect 5940 -460 5950 -399
rect 6010 -460 6020 -399
rect 5940 -470 6020 -460
rect 6990 -400 7070 -310
rect 6990 -460 7000 -400
rect 7060 -460 7070 -400
rect 6990 -470 7070 -460
rect 7120 -400 7200 -140
rect 8310 -100 8320 -40
rect 8380 -100 8390 -40
rect 8310 -230 8390 -100
rect 8310 -290 8320 -230
rect 8380 -290 8390 -230
rect 8310 -300 8390 -290
rect 8520 -190 8600 -180
rect 8520 -250 8530 -190
rect 8590 -250 8600 -190
rect 7120 -460 7130 -400
rect 7190 -460 7200 -400
rect 7120 -470 7200 -460
rect 7260 -400 7340 -390
rect 7260 -460 7270 -400
rect 7330 -460 7340 -400
rect 7260 -470 7340 -460
rect 8520 -400 8600 -250
rect 8650 -190 8730 370
rect 9050 260 9130 410
rect 9440 340 9520 350
rect 9440 280 9450 340
rect 9510 280 9520 340
rect 9050 200 9060 260
rect 9120 200 9130 260
rect 9050 190 9130 200
rect 9210 260 9310 280
rect 9440 270 9520 280
rect 9210 200 9220 260
rect 9280 200 9310 260
rect 9210 190 9310 200
rect 9210 160 9290 190
rect 9190 130 9290 160
rect 9190 70 9210 130
rect 9270 70 9290 130
rect 9190 50 9290 70
rect 8650 -250 8660 -190
rect 8720 -250 8730 -190
rect 8650 -260 8730 -250
rect 8520 -460 8530 -400
rect 8590 -460 8600 -400
rect 8520 -470 8600 -460
rect 8780 -330 8860 -320
rect 8780 -390 8790 -330
rect 8850 -390 8860 -330
rect 8780 -410 8860 -390
rect 8780 -470 8790 -410
rect 8850 -470 8860 -410
rect 8780 -480 8860 -470
rect 8670 -510 8750 -500
rect 6780 -520 6860 -510
rect 6780 -610 6790 -520
rect 6850 -610 6860 -520
rect 8370 -550 8450 -540
rect 8370 -610 8380 -550
rect 8440 -610 8450 -550
rect 8670 -570 8680 -510
rect 8740 -570 8750 -510
rect 8670 -580 8750 -570
rect 5800 -720 5810 -660
rect 5870 -720 5880 -660
rect 5800 -730 5880 -720
rect 5670 -930 5680 -870
rect 5740 -930 5750 -870
rect 6360 -900 6460 -880
rect 5670 -940 5750 -930
rect 6030 -910 6460 -900
rect 6030 -970 6050 -910
rect 6110 -970 6390 -910
rect 6450 -970 6460 -910
rect 6030 -980 6460 -970
rect 6850 -910 6930 -900
rect 6850 -970 6860 -910
rect 6920 -970 6930 -910
rect 5540 -1140 5550 -1080
rect 5610 -1140 5620 -1080
rect 5670 -1070 5750 -1060
rect 5670 -1130 5680 -1070
rect 5740 -1130 5750 -1070
rect 5670 -1140 5750 -1130
rect 6850 -1080 6930 -970
rect 8370 -1010 8450 -610
rect 8370 -1070 8380 -1010
rect 8440 -1070 8450 -1010
rect 8870 -1000 9120 -990
rect 8870 -1060 8880 -1000
rect 8940 -1060 9050 -1000
rect 9110 -1060 9120 -1000
rect 6850 -1140 6860 -1080
rect 6920 -1140 6930 -1080
rect 5540 -1150 5620 -1140
rect 6850 -1150 6930 -1140
rect 6970 -1080 7050 -1070
rect 8370 -1080 8450 -1070
rect 8490 -1070 8570 -1060
rect 8870 -1070 9120 -1060
rect 6970 -1140 6980 -1080
rect 7040 -1140 7050 -1080
rect 8490 -1130 8500 -1070
rect 8560 -1130 8570 -1070
rect 8490 -1140 8570 -1130
rect 6970 -1150 7050 -1140
rect 7280 -1170 7800 -1160
rect 4010 -1220 4110 -1210
rect 1290 -1240 1370 -1220
rect 1290 -1250 1390 -1240
rect 1290 -1330 1300 -1250
rect 1380 -1330 1390 -1250
rect 4010 -1300 4020 -1220
rect 4100 -1300 4110 -1220
rect 7280 -1230 7290 -1170
rect 7350 -1230 7730 -1170
rect 7790 -1230 7800 -1170
rect 7280 -1240 7800 -1230
rect 4010 -1310 4110 -1300
rect 1290 -1340 1390 -1330
<< via2 >>
rect 20 380 80 440
rect 660 380 720 440
rect 190 100 250 160
rect 1210 380 1270 440
rect 1910 370 1970 430
rect 2690 440 2750 500
rect 2280 280 2340 340
rect 3420 440 3480 500
rect 560 100 620 160
rect 1410 90 1470 150
rect 190 -50 250 10
rect 370 -50 430 10
rect 30 -280 90 -220
rect 1430 -120 1490 -60
rect 470 -460 530 -400
rect 2020 80 2080 141
rect 3050 260 3130 270
rect 3050 200 3060 260
rect 3060 200 3120 260
rect 3120 200 3130 260
rect 3050 190 3130 200
rect 3970 370 4030 430
rect 4730 360 4790 420
rect 5510 400 5570 460
rect 5080 290 5140 349
rect 6220 390 6280 450
rect 2860 40 2920 100
rect 3290 40 3350 100
rect 4170 60 4230 121
rect 1600 -120 1660 -60
rect 4180 -90 4240 -30
rect 1560 -270 1620 -210
rect 2830 -310 2910 -230
rect 3990 -280 4050 -220
rect 1690 -460 1750 -400
rect 3130 -400 3210 -390
rect 3130 -460 3140 -400
rect 3140 -460 3200 -400
rect 3200 -460 3210 -400
rect 3130 -470 3210 -460
rect 5870 250 5930 310
rect 6790 390 6850 450
rect 6590 290 6650 350
rect 7530 380 7590 440
rect 8300 440 8360 500
rect 4840 60 4900 119
rect 5690 60 5750 120
rect 6370 40 6430 100
rect 7180 190 7240 250
rect 7910 270 7970 330
rect 9040 420 9120 500
rect 6990 30 7050 90
rect 7410 40 7470 100
rect 8500 70 8560 130
rect 4370 -90 4430 -30
rect 7130 -140 7190 -80
rect 5810 -280 5870 -220
rect 4450 -460 4510 -400
rect 400 -580 450 -570
rect 450 -580 460 -570
rect 400 -630 460 -580
rect 1230 -580 1290 -560
rect 1230 -620 1290 -580
rect 3040 -580 3100 -560
rect 3040 -620 3100 -580
rect 2660 -770 2720 -710
rect 4340 -770 4400 -710
rect 70 -1010 130 -950
rect 2730 -980 2810 -900
rect 190 -1130 250 -1120
rect 190 -1180 250 -1130
rect 1400 -1080 1480 -1070
rect 1400 -1140 1410 -1080
rect 1410 -1140 1470 -1080
rect 1470 -1140 1480 -1080
rect 1400 -1150 1480 -1140
rect 2840 -1070 2920 -1060
rect 2840 -1130 2850 -1070
rect 2850 -1130 2910 -1070
rect 2910 -1130 2920 -1070
rect 2840 -1140 2920 -1130
rect 5550 -720 5610 -660
rect 3620 -1130 3680 -1070
rect 4770 -1060 4830 -1000
rect 7000 -310 7060 -250
rect 5950 -460 6010 -400
rect 8320 -100 8380 -40
rect 8530 -250 8590 -190
rect 7270 -460 7330 -400
rect 9450 280 9510 340
rect 9210 70 9270 130
rect 8660 -250 8720 -190
rect 8790 -390 8850 -330
rect 6790 -580 6850 -550
rect 6790 -610 6850 -580
rect 8380 -610 8440 -550
rect 8680 -570 8740 -510
rect 5810 -720 5870 -660
rect 5680 -930 5740 -870
rect 6390 -970 6450 -910
rect 6860 -970 6920 -910
rect 5680 -1130 5740 -1070
rect 9050 -1060 9110 -1000
rect 6980 -1140 7040 -1080
rect 8500 -1130 8560 -1070
rect 1300 -1330 1380 -1250
rect 4020 -1300 4100 -1220
rect 7730 -1230 7790 -1170
<< metal3 >>
rect 2670 520 3540 530
rect 0 450 800 460
rect 0 370 10 450
rect 92 440 800 450
rect 92 380 660 440
rect 720 380 800 440
rect 92 370 800 380
rect 0 360 800 370
rect 1190 450 2050 460
rect 1190 370 1200 450
rect 1280 430 2050 450
rect 2670 440 2680 520
rect 2760 500 3540 520
rect 2760 440 3420 500
rect 3480 440 3540 500
rect 8290 500 9170 510
rect 5490 470 6352 480
rect 2670 430 3540 440
rect 3950 440 4140 450
rect 1280 370 1910 430
rect 1970 370 2050 430
rect 1190 360 2050 370
rect 3950 360 3960 440
rect 4040 430 4140 440
rect 4040 420 4820 430
rect 4040 360 4730 420
rect 4790 360 4820 420
rect 5490 390 5500 470
rect 5580 450 6352 470
rect 5580 390 6220 450
rect 6280 390 6352 450
rect 5490 380 6352 390
rect 6780 460 7640 470
rect 6780 380 6790 460
rect 6870 440 7640 460
rect 6870 380 7530 440
rect 7590 380 7640 440
rect 8290 420 8300 500
rect 8380 420 9040 500
rect 9120 420 9170 500
rect 8290 410 8640 420
rect 8750 410 9170 420
rect 6780 370 7640 380
rect 2260 350 2360 360
rect 1030 340 1130 350
rect 1030 260 1040 340
rect 1120 260 1130 340
rect 2260 270 2270 350
rect 2350 270 2360 350
rect 3770 350 3870 360
rect 3950 350 4820 360
rect 5060 360 5160 370
rect 2260 260 2360 270
rect 3040 270 3140 280
rect 1030 250 1130 260
rect 3040 190 3050 270
rect 3130 190 3140 270
rect 3770 270 3780 350
rect 3860 270 3870 350
rect 5060 280 5070 360
rect 5150 280 5160 360
rect 6570 360 6670 370
rect 5060 270 5160 280
rect 5860 310 6030 320
rect 3770 260 3870 270
rect 5860 250 5870 310
rect 5930 250 5940 310
rect 5860 240 5940 250
rect 5930 230 5940 240
rect 6020 230 6030 310
rect 6570 270 6580 360
rect 6660 270 6670 360
rect 9430 350 9530 360
rect 7890 340 7990 350
rect 7890 260 7900 340
rect 7980 260 7990 340
rect 9430 270 9440 350
rect 9520 270 9530 350
rect 9430 260 9530 270
rect 5930 220 6030 230
rect 7170 250 7650 260
rect 7890 250 7990 260
rect 3040 180 3140 190
rect 7170 190 7180 250
rect 7240 190 7560 250
rect 7170 180 7560 190
rect 180 170 680 180
rect 7550 170 7560 180
rect 7640 170 7650 250
rect 180 90 190 170
rect 260 160 680 170
rect 260 100 560 160
rect 620 100 680 160
rect 260 90 680 100
rect 180 80 680 90
rect 1390 160 2140 170
rect 7550 160 7650 170
rect 1390 80 1400 160
rect 1480 141 2140 160
rect 1480 80 2020 141
rect 2080 80 2140 141
rect 8490 140 9320 150
rect 4150 130 4930 140
rect 8570 130 9320 140
rect 1390 70 2140 80
rect 2840 110 3360 120
rect 2840 30 2850 110
rect 2930 100 3360 110
rect 2930 40 3290 100
rect 3350 40 3360 100
rect 4150 50 4160 130
rect 4240 119 4930 130
rect 4240 60 4840 119
rect 4900 60 4930 119
rect 4240 50 4930 60
rect 4150 40 4930 50
rect 5670 120 6450 130
rect 5670 40 5680 120
rect 5760 100 6450 120
rect 5760 40 6370 100
rect 6430 40 6450 100
rect 2930 30 3360 40
rect 5670 30 6450 40
rect 6980 100 7490 120
rect 6980 90 7410 100
rect 6980 30 6990 90
rect 7050 40 7410 90
rect 7470 40 7490 100
rect 8570 70 9210 130
rect 9270 70 9320 130
rect 8570 60 9320 70
rect 8490 50 9320 60
rect 7050 30 7490 40
rect 2840 20 3360 30
rect 6980 20 7490 30
rect 180 10 440 20
rect 180 -50 190 10
rect 250 -50 370 10
rect 430 -50 440 10
rect 9020 -20 9120 -10
rect 4170 -30 4440 -20
rect 9020 -30 9030 -20
rect 180 -60 440 -50
rect 1420 -60 1690 -50
rect 180 -80 280 -60
rect 1420 -120 1430 -60
rect 1490 -120 1600 -60
rect 1660 -120 1690 -60
rect 4170 -90 4180 -30
rect 4240 -90 4370 -30
rect 4430 -90 4440 -30
rect 8310 -40 9030 -30
rect 4170 -100 4440 -90
rect 5580 -80 7430 -70
rect 1420 -130 1690 -120
rect 5580 -140 7130 -80
rect 7190 -140 7340 -80
rect 5580 -150 7340 -140
rect 7330 -160 7340 -150
rect 7420 -160 7430 -80
rect 8310 -100 8320 -40
rect 8380 -100 9030 -40
rect 9110 -30 9120 -20
rect 9110 -100 9340 -30
rect 8310 -110 9340 -100
rect 7330 -170 7430 -160
rect 8520 -190 8780 -180
rect 20 -210 1830 -200
rect 20 -220 1560 -210
rect 20 -280 30 -220
rect 90 -270 1560 -220
rect 1620 -270 1830 -210
rect 3980 -220 5880 -210
rect 90 -280 1830 -270
rect 2820 -230 2920 -220
rect 20 -290 100 -280
rect 2820 -310 2830 -230
rect 2910 -240 2920 -230
rect 3030 -230 3130 -220
rect 3030 -240 3040 -230
rect 2910 -310 3040 -240
rect 3120 -310 3130 -230
rect 3980 -280 3990 -220
rect 4050 -280 5810 -220
rect 5870 -280 5880 -220
rect 7540 -230 7640 -220
rect 7540 -240 7550 -230
rect 3980 -290 5880 -280
rect 6990 -250 7550 -240
rect 2820 -320 3130 -310
rect 6990 -310 7000 -250
rect 7060 -310 7550 -250
rect 7630 -310 7640 -230
rect 8520 -250 8530 -190
rect 8590 -250 8660 -190
rect 8720 -250 8780 -190
rect 8520 -260 8780 -250
rect 6990 -320 7640 -310
rect 9420 -310 9520 -300
rect 9420 -320 9430 -310
rect 8780 -330 9430 -320
rect 2240 -380 2340 -370
rect 3760 -380 3860 -370
rect 2240 -390 2250 -380
rect 450 -400 550 -390
rect 450 -480 460 -400
rect 540 -480 550 -400
rect 1680 -400 2250 -390
rect 1680 -460 1690 -400
rect 1750 -460 2250 -400
rect 2330 -460 2340 -380
rect 1680 -470 2340 -460
rect 3120 -390 3220 -380
rect 3760 -390 3770 -380
rect 3120 -470 3130 -390
rect 3210 -460 3770 -390
rect 3850 -460 3860 -380
rect 5050 -380 5150 -370
rect 5050 -390 5060 -380
rect 3210 -470 3860 -460
rect 4440 -400 5060 -390
rect 4440 -460 4450 -400
rect 4510 -460 5060 -400
rect 5140 -460 5150 -380
rect 6570 -380 6670 -370
rect 6570 -390 6580 -380
rect 4440 -470 5150 -460
rect 5940 -400 6580 -390
rect 5940 -460 5950 -400
rect 6010 -460 6580 -400
rect 6660 -460 6670 -380
rect 7880 -380 7980 -370
rect 7880 -389 7890 -380
rect 7460 -390 7890 -389
rect 5940 -470 6670 -460
rect 7260 -400 7890 -390
rect 7260 -460 7270 -400
rect 7330 -460 7890 -400
rect 7970 -460 7980 -380
rect 8780 -390 8790 -330
rect 8850 -390 9430 -330
rect 9510 -390 9520 -310
rect 8780 -400 9520 -390
rect 7260 -470 7980 -460
rect 3120 -480 3220 -470
rect 450 -500 550 -480
rect 8670 -510 8750 -500
rect 8670 -540 8680 -510
rect 1020 -560 1120 -540
rect 3020 -550 3120 -540
rect 380 -570 1030 -560
rect 380 -630 400 -570
rect 460 -630 1030 -570
rect 380 -640 1030 -630
rect 1110 -640 1120 -560
rect 1220 -560 3030 -550
rect 1220 -620 1230 -560
rect 1290 -620 3030 -560
rect 3110 -620 3120 -550
rect 6780 -550 8680 -540
rect 6780 -610 6790 -550
rect 6850 -610 8380 -550
rect 8440 -570 8680 -550
rect 8740 -570 8750 -510
rect 8440 -610 8750 -570
rect 6780 -620 8750 -610
rect 1220 -630 3120 -620
rect 1020 -650 1120 -640
rect 5540 -660 5880 -650
rect 2650 -710 4410 -700
rect 2650 -770 2660 -710
rect 2720 -770 4340 -710
rect 4400 -770 4410 -710
rect 5540 -720 5550 -660
rect 5610 -720 5810 -660
rect 5870 -720 5880 -660
rect 5540 -730 5880 -720
rect 2650 -780 4410 -770
rect 5920 -850 6020 -840
rect 5920 -860 5930 -850
rect 810 -870 910 -860
rect 450 -930 550 -920
rect 450 -940 460 -930
rect 60 -950 460 -940
rect 60 -1010 70 -950
rect 130 -1010 460 -950
rect 540 -1010 550 -930
rect 810 -950 820 -870
rect 900 -950 910 -870
rect 5670 -870 5930 -860
rect 3760 -890 3860 -880
rect 810 -960 910 -950
rect 2020 -900 2120 -890
rect 820 -990 900 -960
rect 2020 -980 2030 -900
rect 2110 -980 2120 -900
rect 2020 -990 2120 -980
rect 2720 -900 3770 -890
rect 2720 -980 2730 -900
rect 2810 -960 3770 -900
rect 3850 -960 3860 -890
rect 5670 -930 5680 -870
rect 5740 -930 5930 -870
rect 6010 -930 6020 -850
rect 2810 -970 3860 -960
rect 2810 -980 2820 -970
rect 4760 -980 4840 -930
rect 5670 -940 6020 -930
rect 6360 -890 6460 -880
rect 6360 -970 6370 -890
rect 6450 -970 6460 -890
rect 7870 -890 7970 -880
rect 7870 -900 7880 -890
rect 6360 -980 6460 -970
rect 6850 -910 7880 -900
rect 6850 -970 6860 -910
rect 6920 -970 7880 -910
rect 7960 -970 7970 -890
rect 6850 -980 7970 -970
rect 9020 -980 9120 -970
rect 2720 -990 2820 -980
rect 4750 -990 4850 -980
rect 60 -1020 550 -1010
rect 3010 -1050 3110 -1040
rect 1730 -1060 1830 -1050
rect 1390 -1070 1490 -1060
rect 1730 -1070 1740 -1060
rect 1020 -1100 1120 -1090
rect 1020 -1110 1030 -1100
rect 180 -1120 1030 -1110
rect 180 -1180 190 -1120
rect 250 -1180 1030 -1120
rect 1110 -1180 1120 -1100
rect 1390 -1150 1400 -1070
rect 1480 -1140 1740 -1070
rect 1820 -1140 1830 -1060
rect 1480 -1150 1830 -1140
rect 2830 -1060 2930 -1050
rect 3010 -1060 3020 -1050
rect 2830 -1140 2840 -1060
rect 2920 -1130 3020 -1060
rect 3100 -1130 3110 -1050
rect 2920 -1140 3110 -1130
rect 3600 -1060 3700 -1050
rect 3600 -1140 3610 -1060
rect 3690 -1140 3700 -1060
rect 4750 -1070 4760 -990
rect 4840 -1070 4850 -990
rect 6570 -1050 6670 -1040
rect 6570 -1060 6580 -1050
rect 4750 -1080 4850 -1070
rect 5670 -1070 6580 -1060
rect 5670 -1130 5680 -1070
rect 5740 -1130 6580 -1070
rect 6660 -1130 6670 -1050
rect 7330 -1060 7430 -1050
rect 9020 -1060 9030 -980
rect 9110 -1060 9120 -980
rect 9410 -1050 9510 -1040
rect 9410 -1060 9420 -1050
rect 7330 -1070 7340 -1060
rect 5670 -1140 6670 -1130
rect 6970 -1080 7340 -1070
rect 6970 -1140 6980 -1080
rect 7040 -1140 7340 -1080
rect 7420 -1140 7430 -1060
rect 8490 -1070 9420 -1060
rect 8490 -1130 8500 -1070
rect 8560 -1130 9420 -1070
rect 9500 -1130 9510 -1050
rect 8490 -1140 9510 -1130
rect 2830 -1150 2930 -1140
rect 3600 -1150 3700 -1140
rect 6970 -1150 7430 -1140
rect 7700 -1150 7800 -1140
rect 1390 -1160 1490 -1150
rect 180 -1190 1120 -1180
rect 2210 -1210 2330 -1200
rect 1290 -1240 1370 -1220
rect 2210 -1240 2240 -1210
rect 1290 -1250 2240 -1240
rect 1290 -1330 1300 -1250
rect 1380 -1290 2240 -1250
rect 2320 -1290 2330 -1210
rect 3610 -1220 3690 -1150
rect 5050 -1210 5150 -1200
rect 4010 -1220 4110 -1210
rect 5050 -1220 5060 -1210
rect 1380 -1300 2330 -1290
rect 4010 -1300 4020 -1220
rect 4100 -1290 5060 -1220
rect 5140 -1290 5150 -1210
rect 7700 -1230 7710 -1150
rect 7790 -1230 7800 -1150
rect 7700 -1240 7800 -1230
rect 4100 -1300 5150 -1290
rect 1380 -1330 1390 -1300
rect 4010 -1310 4110 -1300
rect 1290 -1340 1390 -1330
<< via3 >>
rect 10 440 92 450
rect 10 380 20 440
rect 20 380 80 440
rect 80 380 92 440
rect 10 370 92 380
rect 1200 440 1280 450
rect 1200 380 1210 440
rect 1210 380 1270 440
rect 1270 380 1280 440
rect 2680 500 2760 520
rect 2680 440 2690 500
rect 2690 440 2750 500
rect 2750 440 2760 500
rect 1200 370 1280 380
rect 3960 430 4040 440
rect 3960 370 3970 430
rect 3970 370 4030 430
rect 4030 370 4040 430
rect 3960 360 4040 370
rect 5500 460 5580 470
rect 5500 400 5510 460
rect 5510 400 5570 460
rect 5570 400 5580 460
rect 5500 390 5580 400
rect 6790 450 6870 460
rect 6790 390 6850 450
rect 6850 390 6870 450
rect 6790 380 6870 390
rect 8300 440 8360 500
rect 8360 440 8380 500
rect 8300 420 8380 440
rect 1040 260 1120 340
rect 2270 340 2350 350
rect 2270 280 2280 340
rect 2280 280 2340 340
rect 2340 280 2350 340
rect 2270 270 2350 280
rect 3050 190 3130 270
rect 3780 270 3860 350
rect 5070 349 5150 360
rect 5070 290 5080 349
rect 5080 290 5140 349
rect 5140 290 5150 349
rect 5070 280 5150 290
rect 5940 230 6020 310
rect 6580 350 6660 360
rect 6580 290 6590 350
rect 6590 290 6650 350
rect 6650 290 6660 350
rect 6580 270 6660 290
rect 7900 330 7980 340
rect 7900 270 7910 330
rect 7910 270 7970 330
rect 7970 270 7980 330
rect 7900 260 7980 270
rect 9440 340 9520 350
rect 9440 280 9450 340
rect 9450 280 9510 340
rect 9510 280 9520 340
rect 9440 270 9520 280
rect 7560 170 7640 250
rect 190 160 260 170
rect 190 100 250 160
rect 250 100 260 160
rect 190 90 260 100
rect 1400 150 1480 160
rect 1400 90 1410 150
rect 1410 90 1470 150
rect 1470 90 1480 150
rect 1400 80 1480 90
rect 8490 130 8570 140
rect 2850 100 2930 110
rect 2850 40 2860 100
rect 2860 40 2920 100
rect 2920 40 2930 100
rect 4160 121 4240 130
rect 4160 60 4170 121
rect 4170 60 4230 121
rect 4230 60 4240 121
rect 4160 50 4240 60
rect 5680 60 5690 120
rect 5690 60 5750 120
rect 5750 60 5760 120
rect 5680 40 5760 60
rect 2850 30 2930 40
rect 8490 70 8500 130
rect 8500 70 8560 130
rect 8560 70 8570 130
rect 8490 60 8570 70
rect 7340 -160 7420 -80
rect 9030 -100 9110 -20
rect 3040 -310 3120 -230
rect 7550 -310 7630 -230
rect 460 -460 470 -400
rect 470 -460 530 -400
rect 530 -460 540 -400
rect 460 -480 540 -460
rect 2250 -460 2330 -380
rect 3770 -460 3850 -380
rect 5060 -460 5140 -380
rect 6580 -460 6660 -380
rect 7890 -460 7970 -380
rect 9430 -390 9510 -310
rect 1030 -640 1110 -560
rect 3030 -560 3110 -550
rect 3030 -620 3040 -560
rect 3040 -620 3100 -560
rect 3100 -620 3110 -560
rect 460 -1010 540 -930
rect 820 -950 900 -870
rect 2030 -980 2110 -900
rect 3770 -960 3850 -890
rect 5930 -930 6010 -850
rect 6370 -910 6450 -890
rect 6370 -970 6390 -910
rect 6390 -970 6450 -910
rect 7880 -970 7960 -890
rect 1030 -1180 1110 -1100
rect 1400 -1150 1480 -1070
rect 1740 -1140 1820 -1060
rect 3020 -1130 3100 -1050
rect 3610 -1070 3690 -1060
rect 3610 -1130 3620 -1070
rect 3620 -1130 3680 -1070
rect 3680 -1130 3690 -1070
rect 3610 -1140 3690 -1130
rect 4760 -1000 4840 -990
rect 4760 -1060 4770 -1000
rect 4770 -1060 4830 -1000
rect 4830 -1060 4840 -1000
rect 4760 -1070 4840 -1060
rect 6580 -1130 6660 -1050
rect 9030 -1000 9110 -980
rect 9030 -1060 9050 -1000
rect 9050 -1060 9110 -1000
rect 7340 -1140 7420 -1060
rect 9420 -1130 9500 -1050
rect 2240 -1290 2320 -1210
rect 5060 -1290 5140 -1210
rect 7710 -1170 7790 -1150
rect 7710 -1230 7730 -1170
rect 7730 -1230 7790 -1170
<< metal4 >>
rect 10 460 90 640
rect 0 450 100 460
rect 0 370 10 450
rect 92 370 100 450
rect 0 360 100 370
rect 190 180 270 630
rect 180 170 270 180
rect 180 90 190 170
rect 260 90 270 170
rect 180 80 270 90
rect 450 -390 540 630
rect 450 -400 550 -390
rect 450 -480 460 -400
rect 540 -480 550 -400
rect 450 -500 550 -480
rect 470 -920 550 -500
rect 820 -860 900 630
rect 1200 460 1280 650
rect 1190 450 1290 460
rect 1190 370 1200 450
rect 1280 370 1290 450
rect 1190 360 1290 370
rect 1030 340 1130 350
rect 1030 260 1040 340
rect 1120 260 1130 340
rect 1030 250 1130 260
rect 1040 -540 1120 250
rect 1400 170 1480 670
rect 1390 160 1490 170
rect 1390 80 1400 160
rect 1480 80 1490 160
rect 1390 70 1490 80
rect 1020 -560 1120 -540
rect 1020 -640 1030 -560
rect 1110 -640 1120 -560
rect 1020 -650 1120 -640
rect 450 -930 550 -920
rect 450 -1010 460 -930
rect 540 -1010 550 -930
rect 810 -870 910 -860
rect 810 -950 820 -870
rect 900 -950 910 -870
rect 810 -960 910 -950
rect 450 -1020 550 -1010
rect 1040 -1020 1120 -650
rect 930 -1100 1120 -1020
rect 1750 -1050 1830 -200
rect 2040 -890 2120 630
rect 2680 530 2760 640
rect 2670 520 2770 530
rect 2670 440 2680 520
rect 2760 440 2770 520
rect 2670 430 2770 440
rect 2260 350 2360 360
rect 2260 270 2270 350
rect 2350 270 2360 350
rect 2260 260 2360 270
rect 2280 -370 2340 260
rect 2850 120 2930 640
rect 3040 270 3140 280
rect 3040 190 3050 270
rect 3130 190 3140 270
rect 3040 180 3140 190
rect 2840 110 2960 120
rect 2840 30 2850 110
rect 2930 30 2960 110
rect 2840 20 2960 30
rect 3050 -220 3130 180
rect 3030 -230 3130 -220
rect 3030 -310 3040 -230
rect 3120 -310 3130 -230
rect 3030 -320 3130 -310
rect 2240 -380 2340 -370
rect 2240 -460 2250 -380
rect 2330 -460 2340 -380
rect 2240 -470 2340 -460
rect 2020 -900 2120 -890
rect 2020 -980 2030 -900
rect 2110 -980 2120 -900
rect 2020 -990 2120 -980
rect 1730 -1060 1830 -1050
rect 930 -1150 1030 -1100
rect 1020 -1180 1030 -1150
rect 1110 -1180 1120 -1100
rect 1390 -1070 1490 -1060
rect 1390 -1150 1400 -1070
rect 1480 -1150 1490 -1070
rect 1730 -1140 1740 -1060
rect 1820 -1140 1830 -1060
rect 1730 -1150 1830 -1140
rect 1390 -1160 1490 -1150
rect 1020 -1190 1120 -1180
rect 2250 -1200 2330 -470
rect 3020 -550 3120 -540
rect 3020 -620 3030 -550
rect 3110 -620 3120 -550
rect 3020 -630 3120 -620
rect 3030 -1040 3110 -630
rect 3610 -990 3690 620
rect 3960 450 4040 640
rect 3950 440 4060 450
rect 3950 360 3960 440
rect 4040 360 4060 440
rect 3770 350 3870 360
rect 3950 350 4060 360
rect 3770 270 3780 350
rect 3860 270 3870 350
rect 3770 260 3870 270
rect 3780 -370 3860 260
rect 4160 140 4240 640
rect 4150 130 4250 140
rect 4150 50 4160 130
rect 4240 50 4250 130
rect 4150 40 4250 50
rect 3760 -380 3860 -370
rect 3760 -460 3770 -380
rect 3850 -460 3860 -380
rect 3760 -470 3860 -460
rect 3780 -880 3860 -470
rect 3760 -890 3860 -880
rect 3760 -960 3770 -890
rect 3850 -960 3860 -890
rect 3760 -970 3860 -960
rect 4760 -980 4840 620
rect 5500 480 5580 640
rect 5490 470 5610 480
rect 5490 390 5500 470
rect 5580 390 5610 470
rect 5490 380 5610 390
rect 5060 360 5160 370
rect 5060 280 5070 360
rect 5150 280 5160 360
rect 5060 270 5160 280
rect 5070 -370 5150 270
rect 5680 130 5760 640
rect 5930 310 6030 320
rect 5930 230 5940 310
rect 6020 230 6030 310
rect 5930 220 6030 230
rect 5670 120 5780 130
rect 5670 40 5680 120
rect 5760 40 5780 120
rect 5670 30 5780 40
rect 5050 -380 5150 -370
rect 5050 -460 5060 -380
rect 5140 -460 5150 -380
rect 5050 -470 5150 -460
rect 4750 -990 4850 -980
rect 3010 -1050 3110 -1040
rect 3010 -1130 3020 -1050
rect 3100 -1130 3110 -1050
rect 3010 -1140 3110 -1130
rect 3600 -1060 3700 -1050
rect 3600 -1140 3610 -1060
rect 3690 -1140 3700 -1060
rect 4750 -1070 4760 -990
rect 4840 -1070 4850 -990
rect 4750 -1080 4850 -1070
rect 3600 -1150 3700 -1140
rect 5070 -1200 5150 -470
rect 5940 -840 6020 220
rect 5920 -850 6020 -840
rect 5920 -930 5930 -850
rect 6010 -930 6020 -850
rect 6380 -880 6460 620
rect 6790 470 6870 670
rect 6780 460 6890 470
rect 6780 380 6790 460
rect 6870 380 6890 460
rect 6780 370 6890 380
rect 6570 360 6670 370
rect 6570 270 6580 360
rect 6660 270 6670 360
rect 6570 260 6670 270
rect 6590 -370 6670 260
rect 6990 120 7070 670
rect 7550 250 7650 260
rect 7550 170 7560 250
rect 7640 170 7650 250
rect 7550 160 7650 170
rect 6980 20 7089 120
rect 7330 -80 7430 -70
rect 7330 -160 7340 -80
rect 7420 -160 7430 -80
rect 7330 -170 7430 -160
rect 6570 -380 6670 -370
rect 6570 -460 6580 -380
rect 6660 -460 6670 -380
rect 6570 -470 6670 -460
rect 5920 -940 6020 -930
rect 6360 -890 6460 -880
rect 6360 -970 6370 -890
rect 6450 -970 6460 -890
rect 6360 -980 6460 -970
rect 6590 -1040 6670 -470
rect 6570 -1050 6670 -1040
rect 7350 -1050 7430 -170
rect 7560 -220 7640 160
rect 7540 -230 7640 -220
rect 7540 -310 7550 -230
rect 7630 -310 7640 -230
rect 7540 -320 7640 -310
rect 6570 -1130 6580 -1050
rect 6660 -1130 6670 -1050
rect 6570 -1140 6670 -1130
rect 7330 -1060 7430 -1050
rect 7330 -1140 7340 -1060
rect 7420 -1140 7430 -1060
rect 7720 -1140 7800 640
rect 8300 510 8380 650
rect 8290 500 8430 510
rect 8290 420 8300 500
rect 8380 420 8430 500
rect 8290 410 8430 420
rect 7890 340 7990 350
rect 7890 260 7900 340
rect 7980 260 7990 340
rect 7890 250 7990 260
rect 7900 -370 7980 250
rect 8490 180 8570 650
rect 8480 140 8580 180
rect 8480 60 8490 140
rect 8570 60 8580 140
rect 8480 50 8580 60
rect 9040 -10 9120 620
rect 9020 -20 9120 -10
rect 9020 -100 9030 -20
rect 9110 -100 9120 -20
rect 9020 -110 9120 -100
rect 9260 -110 9340 620
rect 9430 350 9530 360
rect 9430 270 9440 350
rect 9520 270 9530 350
rect 9430 260 9530 270
rect 7880 -380 7980 -370
rect 7880 -460 7890 -380
rect 7970 -460 7980 -380
rect 7880 -470 7980 -460
rect 7890 -880 7970 -470
rect 7870 -890 7970 -880
rect 7870 -970 7880 -890
rect 7960 -970 7970 -890
rect 9040 -970 9120 -110
rect 9440 -300 9520 260
rect 9420 -310 9520 -300
rect 9420 -390 9430 -310
rect 9510 -390 9520 -310
rect 9420 -400 9520 -390
rect 7870 -980 7970 -970
rect 9020 -980 9120 -970
rect 9020 -1060 9030 -980
rect 9110 -1060 9120 -980
rect 9430 -1040 9510 -400
rect 9020 -1070 9120 -1060
rect 9410 -1050 9510 -1040
rect 9410 -1130 9420 -1050
rect 9500 -1130 9510 -1050
rect 9410 -1140 9510 -1130
rect 7330 -1150 7430 -1140
rect 7700 -1150 7800 -1140
rect 2210 -1210 2330 -1200
rect 2210 -1290 2240 -1210
rect 2320 -1290 2330 -1210
rect 2210 -1300 2330 -1290
rect 5050 -1210 5150 -1200
rect 5050 -1290 5060 -1210
rect 5140 -1290 5150 -1210
rect 7700 -1230 7710 -1150
rect 7790 -1230 7800 -1150
rect 7700 -1240 7800 -1230
rect 5050 -1300 5150 -1290
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_0
timestamp 1691611044
transform 1 0 0 0 1 -672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_1
timestamp 1691611044
transform 1 0 1214 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_2
timestamp 1691611044
transform 1 0 2658 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_3
timestamp 1691611044
transform 1 0 3968 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_4
timestamp 1691611044
transform 1 0 5478 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_5
timestamp 1691611044
transform 1 0 6788 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_6
timestamp 1691611044
transform 1 0 8310 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0
timestamp 1691611044
transform 1 0 0 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_1
timestamp 1691611044
transform 1 0 1214 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_2
timestamp 1691611044
transform 1 0 2658 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_3
timestamp 1691611044
transform 1 0 3968 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_4
timestamp 1691611044
transform 1 0 5478 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_5
timestamp 1691611044
transform 1 0 6788 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_6
timestamp 1691611044
transform 1 0 8310 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0
timestamp 1691611044
transform 1 0 728 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1691611044
transform 1 0 1972 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_2
timestamp 1691611044
transform 1 0 9166 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_0
timestamp 1691611044
transform 1 0 620 0 1 -672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_1
timestamp 1691611044
transform 1 0 1840 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_2
timestamp 1691611044
transform 1 0 3290 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_3
timestamp 1691611044
transform 1 0 4600 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_4
timestamp 1691611044
transform 1 0 6118 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_5
timestamp 1691611044
transform 1 0 7428 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_6
timestamp 1691611044
transform 1 0 8982 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_7
timestamp 1691611044
transform 1 0 3360 0 1 -1342
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_8
timestamp 1691611044
transform 1 0 4688 0 1 -1342
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_9
timestamp 1691611044
transform 1 0 6218 0 1 -1342
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_10
timestamp 1691611044
transform 1 0 7518 0 1 -1342
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1691611044
transform 1 0 2448 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1691611044
transform 1 0 5278 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1691611044
transform 1 0 8100 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1691611044
transform 1 0 2448 0 1 -670
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1691611044
transform 1 0 2448 0 1 -1342
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1691611044
transform 1 0 5278 0 1 -668
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1691611044
transform 1 0 5278 0 1 -1342
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1691611044
transform 1 0 8100 0 1 -668
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1691611044
transform 1 0 8100 0 1 -1342
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0
timestamp 1691611044
transform 1 0 480 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1691611044
transform 1 0 1714 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_2
timestamp 1691611044
transform 1 0 3228 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_3
timestamp 1691611044
transform 1 0 4528 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_4
timestamp 1691611044
transform 1 0 6038 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_5
timestamp 1691611044
transform 1 0 7348 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_6
timestamp 1691611044
transform 1 0 8890 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_7
timestamp 1691611044
transform 1 0 0 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_8
timestamp 1691611044
transform 1 0 1214 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_9
timestamp 1691611044
transform 1 0 2658 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_10
timestamp 1691611044
transform 1 0 3968 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_11
timestamp 1691611044
transform 1 0 5478 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_12
timestamp 1691611044
transform 1 0 6788 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_13
timestamp 1691611044
transform 1 0 8308 0 1 -1342
box -38 -48 682 592
<< end >>
