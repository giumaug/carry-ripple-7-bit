magic
tech sky130A
magscale 1 2
timestamp 1740868184
<< nwell >>
rect -40 260 9580 592
rect 2540 -100 2710 -78
rect 2540 -400 2630 -100
rect 2540 -420 2710 -400
rect 3234 -409 3270 -88
rect 3870 -409 3937 -88
rect 4543 -409 4568 -88
rect 5185 -406 5245 -88
rect 5394 -398 5460 -86
rect 5394 -406 5580 -398
rect 5185 -407 5580 -406
rect 6045 -407 6090 -86
rect 6700 -407 6754 -86
rect 7365 -407 7395 -86
rect 8013 -407 8068 -86
rect 8200 -90 8370 -80
rect 8200 -400 8300 -90
rect 5188 -410 5580 -407
rect 8200 -410 8370 -400
rect 8895 -407 8952 -86
rect 5400 -760 5570 -750
rect 671 -1081 692 -760
rect 1120 -1081 1182 -760
rect 1880 -1081 1940 -760
rect 2360 -1081 2417 -760
rect 2570 -1080 2630 -760
rect 5400 -1080 5450 -760
rect 2570 -1090 2750 -1080
rect 5400 -1090 5570 -1080
rect 6155 -1081 6184 -760
rect 7460 -1081 7484 -760
rect 8224 -1081 8276 -760
rect 8986 -1081 9131 -760
<< pwell >>
rect 1109 -49 1235 60
rect 1665 -48 1720 48
<< locali >>
rect 454 527 502 561
rect 1121 527 1217 561
rect 1665 527 1719 561
rect 2349 527 2453 561
rect 2532 527 2668 561
rect 3115 527 3233 561
rect 3866 527 3973 561
rect 4427 527 4530 561
rect 5170 527 5282 561
rect 5363 527 5481 561
rect 5928 527 6044 561
rect 6675 527 6792 561
rect 7246 527 7352 561
rect 7990 527 8104 561
rect 8184 527 8313 561
rect 8759 527 8894 561
rect 10 280 90 300
rect 10 240 30 280
rect 70 240 90 280
rect 10 220 90 240
rect 2026 249 2101 260
rect 2026 243 2051 249
rect 2085 243 2101 249
rect 437 -17 504 17
rect 1117 -17 1221 17
rect 1656 -18 1720 17
rect 2348 -17 2457 17
rect 2526 -17 2661 17
rect 3115 -17 3235 17
rect 3863 -17 3973 17
rect 4417 -17 4534 17
rect 5170 -17 5285 17
rect 5359 -17 5483 17
rect 5925 -17 6047 17
rect 6678 -17 6794 17
rect 7237 -17 7354 17
rect 7981 -17 8104 17
rect 8178 -17 8315 17
rect 8768 -17 8894 17
rect 5110 -109 5280 -104
rect 529 -145 624 -111
rect 1169 -145 1231 -109
rect 1756 -143 1842 -109
rect 2388 -143 2452 -109
rect 2523 -143 2664 -109
rect 3208 -143 3316 -109
rect 3828 -143 3974 -109
rect 4513 -143 4604 -109
rect 5110 -120 5282 -109
rect 5149 -141 5282 -120
rect 5367 -141 5487 -107
rect 6027 -141 6121 -107
rect 6655 -141 6799 -107
rect 7337 -141 7433 -107
rect 7977 -141 8103 -107
rect 8183 -141 8314 -107
rect 8857 -141 8987 -107
rect 545 -689 624 -655
rect 1155 -660 1220 -650
rect 5126 -653 5281 -651
rect 1163 -687 1217 -660
rect 1762 -687 1843 -653
rect 2383 -687 2453 -653
rect 2533 -687 2665 -653
rect 3200 -687 3293 -653
rect 3830 -687 3976 -653
rect 4502 -687 4603 -653
rect 5126 -686 5285 -653
rect 5362 -685 5484 -651
rect 6027 -686 6126 -651
rect 6661 -685 6793 -651
rect 7333 -685 7433 -651
rect 7974 -685 8107 -651
rect 8189 -685 8313 -651
rect 8859 -685 8997 -651
rect 5126 -687 5281 -686
rect 626 -815 732 -781
rect 1092 -815 1222 -781
rect 1844 -815 1977 -781
rect 2332 -815 2451 -781
rect 2537 -815 2660 -781
rect 3293 -815 3364 -781
rect 3895 -815 3973 -781
rect 4600 -815 4692 -781
rect 5233 -815 5283 -781
rect 5369 -815 5490 -781
rect 6111 -815 6226 -781
rect 6763 -815 6792 -781
rect 7425 -815 7523 -781
rect 8060 -815 8106 -781
rect 8187 -815 8318 -781
rect 8944 -815 9174 -781
rect 632 -1359 732 -1325
rect 1087 -1359 1224 -1325
rect 1851 -1359 1975 -1325
rect 2330 -1359 2455 -1325
rect 2528 -1359 2666 -1325
rect 3293 -1359 3363 -1325
rect 3902 -1360 3974 -1325
rect 4603 -1359 4694 -1325
rect 5228 -1359 5285 -1325
rect 5368 -1359 5484 -1325
rect 6113 -1359 6225 -1325
rect 6758 -1359 6811 -1325
rect 7426 -1359 7524 -1325
rect 8062 -1359 8110 -1325
rect 8186 -1359 8313 -1325
rect 8945 -1359 9174 -1325
<< viali >>
rect 30 240 70 280
rect 571 270 606 306
rect 210 220 250 260
rect 680 218 716 253
rect 1240 230 1280 270
rect 1429 215 1463 249
rect 1915 215 1950 251
rect 2051 215 2085 249
rect 2690 220 2730 260
rect 2873 223 2907 258
rect 3320 215 3356 250
rect 3430 210 3470 250
rect 3990 220 4030 260
rect 4181 221 4215 255
rect 4720 210 4760 250
rect 4865 218 4899 253
rect 5507 223 5541 258
rect 5690 220 5730 260
rect 6240 215 6274 249
rect 6375 215 6409 249
rect 6803 225 6840 260
rect 7001 221 7035 255
rect 7433 215 7467 249
rect 7550 217 7584 252
rect 8339 221 8373 255
rect 8525 215 8559 249
rect 9092 215 9126 249
rect 9220 210 9260 250
rect 480 -457 514 -423
rect 390 -570 430 -530
rect 85 -1127 119 -1093
rect 202 -1127 242 -1087
<< metal1 >>
rect 444 496 498 592
rect 1115 496 1218 592
rect 1669 496 1720 592
rect 2354 496 2456 592
rect 2537 496 2661 592
rect 3110 496 3238 592
rect 3851 496 3977 592
rect 4423 496 4532 592
rect 5167 496 5282 592
rect 5367 496 5484 592
rect 5934 496 6044 592
rect 6679 496 6791 592
rect 7240 496 7354 592
rect 7987 496 8105 592
rect 8188 496 8312 592
rect 8765 496 8898 592
rect 550 306 619 330
rect 10 290 90 300
rect 10 230 20 290
rect 80 230 90 290
rect 10 220 90 230
rect 190 260 270 290
rect 550 270 571 306
rect 606 270 619 306
rect 8290 290 8380 310
rect 660 280 740 290
rect 660 270 670 280
rect 550 260 619 270
rect 190 220 210 260
rect 250 220 270 260
rect 190 210 270 220
rect 650 220 670 270
rect 730 270 740 280
rect 1200 280 1310 290
rect 5490 280 5570 290
rect 730 220 760 270
rect 650 218 680 220
rect 716 218 760 220
rect 650 210 760 218
rect 1200 220 1210 280
rect 1270 270 1310 280
rect 1900 270 1980 280
rect 1280 230 1310 270
rect 1270 220 1310 230
rect 1200 210 1310 220
rect 1413 249 1490 270
rect 1413 215 1429 249
rect 1463 215 1490 249
rect 1413 190 1490 215
rect 1900 210 1910 270
rect 1970 210 1980 270
rect 2680 270 2760 280
rect 2026 250 2100 258
rect 1900 200 1980 210
rect 2020 249 2100 250
rect 2020 240 2051 249
rect 2085 240 2100 249
rect 2020 180 2030 240
rect 2090 180 2100 240
rect 2680 210 2690 270
rect 2750 210 2760 270
rect 2680 200 2760 210
rect 2850 270 2930 280
rect 3410 270 3490 280
rect 2850 210 2860 270
rect 2920 210 2930 270
rect 3313 260 3362 270
rect 2850 190 2930 210
rect 3280 250 3362 260
rect 3280 215 3320 250
rect 3356 215 3362 250
rect 3280 199 3362 215
rect 3410 210 3420 270
rect 3480 210 3490 270
rect 3410 200 3490 210
rect 3960 270 4040 280
rect 3960 210 3970 270
rect 4030 210 4040 270
rect 4167 260 4235 265
rect 3960 200 4040 210
rect 4160 255 4240 260
rect 4160 250 4181 255
rect 4215 250 4240 255
rect 3280 190 3360 199
rect 4160 190 4170 250
rect 4230 190 4240 250
rect 4700 210 4720 270
rect 4780 210 4800 270
rect 4700 200 4800 210
rect 4840 260 4920 271
rect 4160 180 4240 190
rect 4840 199 4850 260
rect 4910 199 4920 260
rect 5490 220 5500 280
rect 5560 220 5570 280
rect 5490 210 5570 220
rect 5670 270 5760 280
rect 7520 270 7600 280
rect 5670 210 5680 270
rect 5740 210 5760 270
rect 6780 260 6860 270
rect 2020 170 2100 180
rect 4840 179 4920 199
rect 5670 170 5760 210
rect 6200 250 6330 260
rect 6200 190 6220 250
rect 6280 190 6330 250
rect 6200 170 6330 190
rect 6360 250 6440 260
rect 6360 190 6370 250
rect 6430 190 6440 250
rect 6780 200 6790 260
rect 6850 200 6860 260
rect 6780 190 6860 200
rect 6980 260 7060 270
rect 7520 260 7530 270
rect 6980 200 6990 260
rect 7050 200 7060 260
rect 6980 190 7060 200
rect 7399 250 7480 260
rect 7399 190 7410 250
rect 7470 190 7480 250
rect 7510 210 7530 260
rect 7590 260 7600 270
rect 7590 210 7630 260
rect 8290 230 8300 290
rect 8360 270 8380 290
rect 8360 255 8399 270
rect 8290 221 8339 230
rect 8373 221 8399 255
rect 8290 210 8399 221
rect 8500 260 8590 270
rect 7520 200 7600 210
rect 8500 200 8510 260
rect 8570 200 8590 260
rect 8500 190 8590 200
rect 9050 260 9180 270
rect 9050 200 9060 260
rect 9120 249 9180 260
rect 9126 215 9180 249
rect 9120 200 9180 215
rect 9050 190 9180 200
rect 9210 260 9310 280
rect 9210 200 9220 260
rect 9280 200 9310 260
rect 9210 190 9310 200
rect 6360 180 6440 190
rect 7399 170 7480 190
rect 447 -49 518 48
rect 1114 -49 1223 48
rect 1665 -48 1720 48
rect 2352 17 2461 48
rect 2348 -17 2461 17
rect 2352 -49 2461 -17
rect 2535 -48 2666 48
rect 3111 -48 3238 48
rect 3867 -48 3973 48
rect 4423 -14 4532 48
rect 4422 -48 4651 -14
rect 5166 -48 5285 48
rect 5365 -48 5486 48
rect 5933 -48 6045 48
rect 6675 -48 6794 48
rect 7244 -48 7357 48
rect 7986 -48 8108 48
rect 8185 -48 8314 48
rect 8761 -48 8894 48
rect 541 -176 635 -80
rect 1154 -174 1219 -80
rect 1762 -174 1846 -78
rect 2381 -174 2454 -78
rect 2532 -174 2664 -78
rect 3200 -174 3300 -78
rect 3835 -174 3976 -78
rect 4504 -174 4606 -78
rect 5144 -172 5283 -78
rect 5361 -172 5487 -76
rect 6023 -172 6124 -76
rect 6665 -172 6794 -76
rect 7334 -172 7431 -76
rect 7974 -172 8104 -76
rect 8186 -172 8313 -76
rect 8845 -172 8988 -76
rect 470 -423 550 -390
rect 470 -457 480 -423
rect 514 -457 550 -423
rect 470 -470 550 -457
rect 380 -520 460 -510
rect 380 -580 390 -520
rect 450 -580 460 -520
rect 380 -590 460 -580
rect 537 -720 623 -624
rect 1167 -718 1217 -624
rect 1755 -718 1843 -622
rect 2386 -718 2453 -622
rect 2535 -718 2666 -622
rect 3204 -718 3295 -622
rect 3834 -718 3976 -622
rect 4515 -718 4604 -622
rect 5144 -720 5283 -620
rect 5365 -716 5487 -620
rect 6024 -716 6125 -620
rect 6666 -716 6795 -620
rect 7336 -716 7436 -620
rect 7977 -716 8107 -620
rect 8186 -716 8315 -620
rect 8856 -716 8992 -620
rect 634 -846 735 -750
rect 1086 -846 1219 -750
rect 1851 -846 1983 -750
rect 2335 -846 2454 -750
rect 2535 -846 2662 -750
rect 3298 -846 3364 -750
rect 3902 -846 3974 -750
rect 4606 -846 4693 -750
rect 5232 -846 5284 -750
rect 5366 -846 5484 -750
rect 6116 -846 6225 -750
rect 6756 -846 6806 -750
rect 7424 -846 7523 -750
rect 8065 -846 8112 -750
rect 8181 -846 8314 -750
rect 8937 -846 9175 -750
rect 180 -1070 260 -1060
rect 59 -1080 140 -1070
rect 59 -1140 70 -1080
rect 130 -1140 140 -1080
rect 180 -1130 190 -1070
rect 250 -1130 260 -1070
rect 180 -1140 260 -1130
rect 59 -1150 140 -1140
rect 637 -1390 734 -1294
rect 1090 -1390 1222 -1294
rect 1854 -1390 1980 -1294
rect 2336 -1390 2454 -1294
rect 2534 -1390 2665 -1294
rect 3297 -1390 3364 -1294
rect 3906 -1390 3978 -1294
rect 4606 -1390 4696 -1294
rect 5233 -1390 5292 -1294
rect 5364 -1390 5488 -1294
rect 6116 -1390 6226 -1294
rect 6765 -1390 6813 -1294
rect 7425 -1390 7527 -1294
rect 8065 -1390 8105 -1294
rect 8188 -1390 8316 -1294
rect 8944 -1390 9170 -1294
<< via1 >>
rect 20 280 80 290
rect 20 240 30 280
rect 30 240 70 280
rect 70 240 80 280
rect 20 230 80 240
rect 670 253 730 280
rect 670 220 680 253
rect 680 220 716 253
rect 716 220 730 253
rect 1210 270 1270 280
rect 1210 230 1240 270
rect 1240 230 1270 270
rect 1210 220 1270 230
rect 1910 251 1970 270
rect 1910 215 1915 251
rect 1915 215 1950 251
rect 1950 215 1970 251
rect 1910 210 1970 215
rect 2030 215 2051 240
rect 2051 215 2085 240
rect 2085 215 2090 240
rect 2030 180 2090 215
rect 2690 260 2750 270
rect 2690 220 2730 260
rect 2730 220 2750 260
rect 2690 210 2750 220
rect 2860 258 2920 270
rect 2860 223 2873 258
rect 2873 223 2907 258
rect 2907 223 2920 258
rect 2860 210 2920 223
rect 3420 250 3480 270
rect 3420 210 3430 250
rect 3430 210 3470 250
rect 3470 210 3480 250
rect 3970 260 4030 270
rect 3970 220 3990 260
rect 3990 220 4030 260
rect 3970 210 4030 220
rect 4170 221 4181 250
rect 4181 221 4215 250
rect 4215 221 4230 250
rect 4170 190 4230 221
rect 4720 250 4780 270
rect 4720 210 4760 250
rect 4760 210 4780 250
rect 4850 253 4910 260
rect 4850 218 4865 253
rect 4865 218 4899 253
rect 4899 218 4910 253
rect 4850 199 4910 218
rect 5500 258 5560 280
rect 5500 223 5507 258
rect 5507 223 5541 258
rect 5541 223 5560 258
rect 5500 220 5560 223
rect 5680 260 5740 270
rect 5680 220 5690 260
rect 5690 220 5730 260
rect 5730 220 5740 260
rect 5680 210 5740 220
rect 6220 249 6280 250
rect 6220 215 6240 249
rect 6240 215 6274 249
rect 6274 215 6280 249
rect 6220 190 6280 215
rect 6370 249 6430 250
rect 6370 215 6375 249
rect 6375 215 6409 249
rect 6409 215 6430 249
rect 6370 190 6430 215
rect 6790 225 6803 260
rect 6803 225 6840 260
rect 6840 225 6850 260
rect 6790 200 6850 225
rect 6990 255 7050 260
rect 6990 221 7001 255
rect 7001 221 7035 255
rect 7035 221 7050 255
rect 6990 200 7050 221
rect 7410 249 7470 250
rect 7410 215 7433 249
rect 7433 215 7467 249
rect 7467 215 7470 249
rect 7410 190 7470 215
rect 7530 252 7590 270
rect 7530 217 7550 252
rect 7550 217 7584 252
rect 7584 217 7590 252
rect 7530 210 7590 217
rect 8300 255 8360 290
rect 8300 230 8339 255
rect 8339 230 8360 255
rect 8510 249 8570 260
rect 8510 215 8525 249
rect 8525 215 8559 249
rect 8559 215 8570 249
rect 8510 200 8570 215
rect 9060 249 9120 260
rect 9060 215 9092 249
rect 9092 215 9120 249
rect 9060 200 9120 215
rect 9220 250 9280 260
rect 9220 210 9260 250
rect 9260 210 9280 250
rect 9220 200 9280 210
rect 390 -530 450 -520
rect 390 -570 430 -530
rect 430 -570 450 -530
rect 390 -580 450 -570
rect 70 -1093 130 -1080
rect 70 -1127 85 -1093
rect 85 -1127 119 -1093
rect 119 -1127 130 -1093
rect 70 -1140 130 -1127
rect 190 -1087 250 -1070
rect 190 -1127 202 -1087
rect 202 -1127 242 -1087
rect 242 -1127 250 -1087
rect 190 -1130 250 -1127
<< metal2 >>
rect 2680 500 2760 530
rect 0 440 100 460
rect 0 380 20 440
rect 80 380 100 440
rect 0 360 100 380
rect 660 440 740 460
rect 720 380 740 440
rect 10 290 90 360
rect 10 230 20 290
rect 80 230 90 290
rect 10 220 90 230
rect 190 180 270 290
rect 550 180 630 330
rect 660 280 740 380
rect 1190 440 1280 460
rect 1190 380 1210 440
rect 1270 380 1280 440
rect 1190 360 1280 380
rect 660 220 670 280
rect 730 220 740 280
rect 660 210 740 220
rect 1200 280 1280 360
rect 1900 430 1990 460
rect 1900 370 1910 430
rect 1970 370 1990 430
rect 1900 290 1990 370
rect 1200 220 1210 280
rect 1270 220 1280 280
rect 1890 270 1990 290
rect 1200 210 1280 220
rect 180 160 270 180
rect 180 100 190 160
rect 250 100 270 160
rect 180 80 270 100
rect 540 160 630 180
rect 1413 170 1490 270
rect 1890 210 1910 270
rect 1970 210 1990 270
rect 2680 440 2690 500
rect 2750 440 2760 500
rect 2680 270 2760 440
rect 3410 500 3490 530
rect 3410 440 3420 500
rect 3480 440 3490 500
rect 8290 500 8380 510
rect 5490 460 5570 480
rect 1890 190 1990 210
rect 2020 240 2100 250
rect 540 100 560 160
rect 620 100 630 160
rect 540 80 630 100
rect 1390 150 1490 170
rect 1390 90 1410 150
rect 1470 90 1490 150
rect 1390 70 1490 90
rect 2020 180 2030 240
rect 2090 180 2100 240
rect 2680 210 2690 270
rect 2750 210 2760 270
rect 2680 200 2760 210
rect 2850 270 2930 279
rect 2850 210 2860 270
rect 2920 210 2930 270
rect 3410 270 3490 440
rect 2020 141 2100 180
rect 2080 80 2100 141
rect 2020 69 2100 80
rect 2850 100 2930 210
rect 2850 40 2860 100
rect 2920 40 2930 100
rect 2850 20 2930 40
rect 3280 100 3360 260
rect 3410 210 3420 270
rect 3480 210 3490 270
rect 3410 200 3490 210
rect 3960 430 4040 450
rect 3960 370 3970 430
rect 4030 370 4040 430
rect 3960 270 4040 370
rect 4720 420 4800 430
rect 4720 360 4730 420
rect 4790 360 4800 420
rect 4720 270 4800 360
rect 3960 210 3970 270
rect 4030 210 4040 270
rect 3960 200 4040 210
rect 4160 250 4240 260
rect 3280 40 3290 100
rect 3350 40 3360 100
rect 3280 20 3360 40
rect 4160 190 4170 250
rect 4230 211 4240 250
rect 4230 190 4241 211
rect 4700 210 4720 270
rect 4780 210 4800 270
rect 5490 400 5510 460
rect 5490 280 5570 400
rect 6150 450 6300 480
rect 6150 390 6220 450
rect 6280 390 6300 450
rect 6150 370 6300 390
rect 4700 200 4800 210
rect 4839 260 4920 269
rect 4160 121 4241 190
rect 4839 199 4850 260
rect 4910 199 4920 260
rect 5490 220 5500 280
rect 5560 220 5570 280
rect 5490 210 5570 220
rect 5670 270 5750 280
rect 5670 210 5680 270
rect 5740 210 5750 270
rect 6220 260 6300 370
rect 6780 450 6860 470
rect 6780 390 6790 450
rect 6850 390 6860 450
rect 6780 260 6860 390
rect 7520 440 7600 470
rect 7520 380 7530 440
rect 7590 380 7600 440
rect 7520 270 7600 380
rect 4839 140 4920 199
rect 4160 60 4170 121
rect 4230 60 4241 121
rect 4160 39 4241 60
rect 4810 119 4920 140
rect 4810 60 4840 119
rect 4900 60 4920 119
rect 4810 40 4920 60
rect 5670 130 5750 210
rect 6190 250 6330 260
rect 6190 190 6220 250
rect 6280 190 6330 250
rect 6190 170 6330 190
rect 6360 250 6440 260
rect 6360 190 6370 250
rect 6430 190 6440 250
rect 6780 200 6790 260
rect 6850 200 6860 260
rect 6780 190 6860 200
rect 6980 260 7059 270
rect 6980 200 6990 260
rect 7050 200 7059 260
rect 6360 130 6440 190
rect 5670 120 5790 130
rect 5670 60 5690 120
rect 5750 60 5790 120
rect 4810 39 4840 40
rect 5670 30 5790 60
rect 6339 100 6440 130
rect 6339 40 6370 100
rect 6430 40 6440 100
rect 6339 30 6440 40
rect 6980 90 7059 200
rect 7399 250 7480 260
rect 7399 190 7410 250
rect 7470 190 7480 250
rect 7520 210 7530 270
rect 7590 210 7600 270
rect 8290 440 8300 500
rect 8360 440 8380 500
rect 8290 290 8380 440
rect 9030 500 9130 510
rect 9030 420 9040 500
rect 9120 420 9130 500
rect 9030 410 9130 420
rect 8290 230 8300 290
rect 8360 230 8380 290
rect 8290 210 8380 230
rect 8500 260 8580 270
rect 7520 200 7600 210
rect 8500 200 8510 260
rect 8570 200 8580 260
rect 7399 170 7480 190
rect 8500 180 8580 200
rect 9050 260 9130 410
rect 9050 200 9060 260
rect 9120 200 9130 260
rect 9050 190 9130 200
rect 9210 260 9310 280
rect 9210 200 9220 260
rect 9280 200 9310 260
rect 9210 190 9310 200
rect 7400 120 7480 170
rect 8480 130 8580 180
rect 9210 160 9290 190
rect 6980 30 6990 90
rect 7050 30 7059 90
rect 6980 20 7059 30
rect 7380 100 7490 120
rect 7380 40 7410 100
rect 7470 40 7490 100
rect 8480 70 8500 130
rect 8560 70 8580 130
rect 8480 50 8580 70
rect 9190 130 9290 160
rect 9190 70 9210 130
rect 9270 70 9290 130
rect 9190 50 9290 70
rect 7380 20 7490 40
rect 470 -400 550 -390
rect 530 -460 550 -400
rect 470 -470 550 -460
rect 380 -520 470 -510
rect 380 -580 390 -520
rect 450 -570 470 -520
rect 380 -630 400 -580
rect 460 -630 470 -570
rect 380 -640 470 -630
rect 60 -950 140 -940
rect 60 -1010 70 -950
rect 130 -1010 140 -950
rect 60 -1080 140 -1010
rect 60 -1140 70 -1080
rect 130 -1140 140 -1080
rect 60 -1150 140 -1140
rect 180 -1070 260 -1060
rect 180 -1180 190 -1070
rect 250 -1180 260 -1070
rect 180 -1190 260 -1180
<< via2 >>
rect 20 380 80 440
rect 660 380 720 440
rect 1210 380 1270 440
rect 1910 370 1970 430
rect 190 100 250 160
rect 2690 440 2750 500
rect 3420 440 3480 500
rect 560 100 620 160
rect 1410 90 1470 150
rect 2020 80 2080 141
rect 2860 40 2920 100
rect 3970 370 4030 430
rect 4730 360 4790 420
rect 3290 40 3350 100
rect 5510 400 5570 460
rect 6220 390 6280 450
rect 6790 390 6850 450
rect 7530 380 7590 440
rect 4170 60 4230 121
rect 4840 60 4900 119
rect 5690 60 5750 120
rect 6370 40 6430 100
rect 8300 440 8360 500
rect 9040 420 9120 500
rect 6990 30 7050 90
rect 7410 40 7470 100
rect 8500 70 8560 130
rect 9210 70 9270 130
rect 470 -460 530 -400
rect 400 -580 450 -570
rect 450 -580 460 -570
rect 400 -630 460 -580
rect 70 -1010 130 -950
rect 190 -1130 250 -1120
rect 190 -1180 250 -1130
<< metal3 >>
rect 2670 520 3540 530
rect 0 450 800 460
rect 0 370 10 450
rect 92 440 800 450
rect 92 380 660 440
rect 720 380 800 440
rect 92 370 800 380
rect 0 360 800 370
rect 1190 450 2050 460
rect 1190 370 1200 450
rect 1280 430 2050 450
rect 2670 440 2680 520
rect 2760 500 3540 520
rect 2760 440 3420 500
rect 3480 440 3540 500
rect 8290 500 9170 510
rect 5490 470 6352 480
rect 2670 430 3540 440
rect 3950 440 4140 450
rect 1280 370 1910 430
rect 1970 370 2050 430
rect 1190 360 2050 370
rect 3950 360 3960 440
rect 4040 430 4140 440
rect 4040 420 4820 430
rect 4040 360 4730 420
rect 4790 360 4820 420
rect 5490 390 5500 470
rect 5580 450 6352 470
rect 5580 390 6220 450
rect 6280 390 6352 450
rect 5490 380 6352 390
rect 6780 460 7640 470
rect 6780 380 6790 460
rect 6870 440 7640 460
rect 6870 380 7530 440
rect 7590 380 7640 440
rect 8290 420 8300 500
rect 8380 420 9040 500
rect 9120 420 9170 500
rect 8290 410 9170 420
rect 6780 370 7640 380
rect 3950 350 4820 360
rect 180 170 680 180
rect 180 90 190 170
rect 260 160 680 170
rect 260 100 560 160
rect 620 100 680 160
rect 260 90 680 100
rect 180 80 680 90
rect 1390 160 2140 170
rect 1390 80 1400 160
rect 1480 141 2140 160
rect 1480 80 2020 141
rect 2080 80 2140 141
rect 8490 140 9320 150
rect 4150 130 4930 140
rect 8570 130 9320 140
rect 1390 70 2140 80
rect 2840 110 3360 120
rect 2840 30 2850 110
rect 2930 100 3360 110
rect 2930 40 3290 100
rect 3350 40 3360 100
rect 4150 50 4160 130
rect 4240 119 4930 130
rect 4240 60 4840 119
rect 4900 60 4930 119
rect 4240 50 4930 60
rect 4150 40 4930 50
rect 5670 120 6450 130
rect 5670 40 5680 120
rect 5760 100 6450 120
rect 5760 40 6370 100
rect 6430 40 6450 100
rect 2930 30 3360 40
rect 5670 30 6450 40
rect 6980 100 7490 120
rect 6980 90 7410 100
rect 6980 30 6990 90
rect 7050 40 7410 90
rect 7470 40 7490 100
rect 8570 70 9210 130
rect 9270 70 9320 130
rect 8570 60 9320 70
rect 8490 50 9320 60
rect 7050 30 7490 40
rect 2840 20 3360 30
rect 6980 20 7490 30
rect 450 -400 550 -390
rect 450 -480 460 -400
rect 540 -480 550 -400
rect 450 -500 550 -480
rect 380 -570 1120 -560
rect 380 -630 400 -570
rect 460 -630 1120 -570
rect 380 -640 1120 -630
rect 450 -930 550 -920
rect 450 -940 460 -930
rect 60 -950 460 -940
rect 60 -1010 70 -950
rect 130 -1010 460 -950
rect 540 -1010 550 -930
rect 60 -1020 550 -1010
rect 1020 -1100 1120 -1090
rect 1020 -1110 1030 -1100
rect 180 -1120 1030 -1110
rect 180 -1180 190 -1120
rect 250 -1180 1030 -1120
rect 1110 -1180 1120 -1100
rect 180 -1190 1120 -1180
<< via3 >>
rect 10 440 92 450
rect 10 380 20 440
rect 20 380 80 440
rect 80 380 92 440
rect 10 370 92 380
rect 1200 440 1280 450
rect 1200 380 1210 440
rect 1210 380 1270 440
rect 1270 380 1280 440
rect 2680 500 2760 520
rect 2680 440 2690 500
rect 2690 440 2750 500
rect 2750 440 2760 500
rect 1200 370 1280 380
rect 3960 430 4040 440
rect 3960 370 3970 430
rect 3970 370 4030 430
rect 4030 370 4040 430
rect 3960 360 4040 370
rect 5500 460 5580 470
rect 5500 400 5510 460
rect 5510 400 5570 460
rect 5570 400 5580 460
rect 5500 390 5580 400
rect 6790 450 6870 460
rect 6790 390 6850 450
rect 6850 390 6870 450
rect 6790 380 6870 390
rect 8300 440 8360 500
rect 8360 440 8380 500
rect 8300 420 8380 440
rect 190 160 260 170
rect 190 100 250 160
rect 250 100 260 160
rect 190 90 260 100
rect 1400 150 1480 160
rect 1400 90 1410 150
rect 1410 90 1470 150
rect 1470 90 1480 150
rect 1400 80 1480 90
rect 8490 130 8570 140
rect 2850 100 2930 110
rect 2850 40 2860 100
rect 2860 40 2920 100
rect 2920 40 2930 100
rect 4160 121 4240 130
rect 4160 60 4170 121
rect 4170 60 4230 121
rect 4230 60 4240 121
rect 4160 50 4240 60
rect 5680 60 5690 120
rect 5690 60 5750 120
rect 5750 60 5760 120
rect 5680 40 5760 60
rect 2850 30 2930 40
rect 8490 70 8500 130
rect 8500 70 8560 130
rect 8560 70 8570 130
rect 8490 60 8570 70
rect 460 -460 470 -400
rect 470 -460 530 -400
rect 530 -460 540 -400
rect 460 -480 540 -460
rect 460 -1010 540 -930
rect 1030 -1180 1110 -1100
<< metal4 >>
rect 10 460 90 640
rect 0 450 100 460
rect 0 370 10 450
rect 92 370 100 450
rect 0 360 100 370
rect 190 180 270 630
rect 180 170 270 180
rect 180 90 190 170
rect 260 90 270 170
rect 180 80 270 90
rect 450 -390 540 630
rect 1200 460 1280 650
rect 1190 450 1290 460
rect 1190 370 1200 450
rect 1280 370 1290 450
rect 1190 360 1290 370
rect 450 -400 550 -390
rect 450 -480 460 -400
rect 540 -480 550 -400
rect 1040 -480 1120 330
rect 1400 170 1480 670
rect 2680 530 2760 640
rect 2670 520 2770 530
rect 2670 440 2680 520
rect 2760 440 2770 520
rect 2670 430 2770 440
rect 1390 160 1490 170
rect 1390 80 1400 160
rect 1480 80 1490 160
rect 2850 120 2930 640
rect 3960 450 4040 640
rect 3950 440 4060 450
rect 3950 360 3960 440
rect 4040 360 4060 440
rect 3950 350 4060 360
rect 4160 140 4240 640
rect 5500 480 5580 640
rect 5490 470 5610 480
rect 5490 390 5500 470
rect 5580 390 5610 470
rect 5490 380 5610 390
rect 4150 130 4350 140
rect 5680 130 5760 640
rect 6790 470 6870 670
rect 6780 460 6890 470
rect 6780 380 6790 460
rect 6870 380 6890 460
rect 6780 370 6890 380
rect 1390 70 1490 80
rect 2840 110 2960 120
rect 2840 30 2850 110
rect 2930 30 2960 110
rect 4150 50 4160 130
rect 4240 50 4350 130
rect 4150 40 4350 50
rect 5670 120 5780 130
rect 6990 120 7070 670
rect 8300 510 8380 650
rect 8290 500 8430 510
rect 8290 420 8300 500
rect 8380 420 8430 500
rect 8290 410 8430 420
rect 8490 180 8570 650
rect 8480 140 8580 180
rect 5670 40 5680 120
rect 5760 40 5780 120
rect 5670 30 5780 40
rect 2840 20 2960 30
rect 6980 20 7089 120
rect 8480 60 8490 140
rect 8570 60 8580 140
rect 8480 50 8580 60
rect 450 -500 550 -480
rect 470 -920 550 -500
rect 1000 -590 1120 -480
rect 450 -930 550 -920
rect 450 -1010 460 -930
rect 540 -1010 550 -930
rect 450 -1020 550 -1010
rect 1040 -1020 1120 -590
rect 930 -1100 1120 -1020
rect 930 -1150 1030 -1100
rect 1020 -1180 1030 -1150
rect 1110 -1180 1120 -1100
rect 1020 -1190 1120 -1180
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_0
timestamp 1691611044
transform 1 0 0 0 1 -672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_1
timestamp 1691611044
transform 1 0 1214 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_2
timestamp 1691611044
transform 1 0 2658 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_3
timestamp 1691611044
transform 1 0 3968 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_4
timestamp 1691611044
transform 1 0 5478 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_5
timestamp 1691611044
transform 1 0 6788 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_6
timestamp 1691611044
transform 1 0 8310 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0
timestamp 1691611044
transform 1 0 0 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_1
timestamp 1691611044
transform 1 0 1214 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_2
timestamp 1691611044
transform 1 0 2658 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_3
timestamp 1691611044
transform 1 0 3968 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_4
timestamp 1691611044
transform 1 0 5478 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_5
timestamp 1691611044
transform 1 0 6788 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_6
timestamp 1691611044
transform 1 0 8310 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0
timestamp 1691611044
transform 1 0 728 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1691611044
transform 1 0 1972 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_2
timestamp 1691611044
transform 1 0 9166 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_0
timestamp 1691611044
transform 1 0 620 0 1 -672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_1
timestamp 1691611044
transform 1 0 1840 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_2
timestamp 1691611044
transform 1 0 3290 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_3
timestamp 1691611044
transform 1 0 4600 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_4
timestamp 1691611044
transform 1 0 6118 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_5
timestamp 1691611044
transform 1 0 7428 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_6
timestamp 1691611044
transform 1 0 8982 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_7
timestamp 1691611044
transform 1 0 3360 0 1 -1342
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_8
timestamp 1691611044
transform 1 0 4688 0 1 -1342
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_9
timestamp 1691611044
transform 1 0 6218 0 1 -1342
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_10
timestamp 1691611044
transform 1 0 7518 0 1 -1342
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1691611044
transform 1 0 2448 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1691611044
transform 1 0 5278 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1691611044
transform 1 0 8100 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1691611044
transform 1 0 2448 0 1 -670
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1691611044
transform 1 0 2448 0 1 -1342
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1691611044
transform 1 0 5278 0 1 -668
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1691611044
transform 1 0 5278 0 1 -1342
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1691611044
transform 1 0 8100 0 1 -668
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1691611044
transform 1 0 8100 0 1 -1342
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0
timestamp 1691611044
transform 1 0 480 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1691611044
transform 1 0 1714 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_2
timestamp 1691611044
transform 1 0 3228 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_3
timestamp 1691611044
transform 1 0 4528 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_4
timestamp 1691611044
transform 1 0 6038 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_5
timestamp 1691611044
transform 1 0 7348 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_6
timestamp 1691611044
transform 1 0 8890 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_7
timestamp 1691611044
transform 1 0 0 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_8
timestamp 1691611044
transform 1 0 1214 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_9
timestamp 1691611044
transform 1 0 2658 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_10
timestamp 1691611044
transform 1 0 3968 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_11
timestamp 1691611044
transform 1 0 5478 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_12
timestamp 1691611044
transform 1 0 6788 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_13
timestamp 1691611044
transform 1 0 8308 0 1 -1342
box -38 -48 682 592
<< end >>
