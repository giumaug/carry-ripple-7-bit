magic
tech sky130A
timestamp 1742991778
<< metal3 >>
rect 2710 22430 14720 22435
rect 2710 22390 2715 22430
rect 2755 22390 3065 22430
rect 3105 22390 3340 22430
rect 3380 22390 3615 22430
rect 3655 22390 3890 22430
rect 3930 22390 4165 22430
rect 4205 22390 4440 22430
rect 4480 22390 4715 22430
rect 4755 22390 4990 22430
rect 5030 22390 14720 22430
rect 2710 22385 14720 22390
rect 3060 22295 14720 22345
rect 3060 22205 14720 22255
rect 3060 22115 14720 22165
rect 3060 22025 14720 22075
rect 400 21980 2760 21985
rect 400 21940 405 21980
rect 445 21940 470 21980
rect 510 21940 535 21980
rect 575 21940 2715 21980
rect 2755 21940 2760 21980
rect 400 21935 2760 21940
rect 3060 21935 14720 21985
rect 3060 21845 14720 21895
rect 3060 21755 14720 21805
rect 3060 21670 14720 21715
rect 3060 21665 14385 21670
rect 3060 21575 14720 21625
rect 3060 21485 14720 21535
rect 3060 21395 14720 21445
rect 3060 21305 14720 21355
rect 3060 21215 14720 21265
rect 3060 21135 14720 21175
rect 3060 21055 14720 21095
rect 3060 20975 14720 21015
rect 3060 20895 14720 20935
rect 3060 20815 14720 20855
rect 3060 20735 14720 20775
rect 3060 20655 14720 20695
rect 3060 20575 14720 20615
rect 3060 20495 14720 20535
<< via3 >>
rect 2715 22390 2755 22430
rect 3065 22390 3105 22430
rect 3340 22390 3380 22430
rect 3615 22390 3655 22430
rect 3890 22390 3930 22430
rect 4165 22390 4205 22430
rect 4440 22390 4480 22430
rect 4715 22390 4755 22430
rect 4990 22390 5030 22430
rect 405 21940 445 21980
rect 470 21940 510 21980
rect 535 21940 575 21980
rect 2715 21940 2755 21980
<< metal4 >>
rect 3067 22485 3097 22576
rect 3343 22485 3373 22576
rect 3619 22485 3649 22576
rect 3895 22485 3925 22576
rect 4171 22485 4201 22576
rect 4447 22485 4477 22576
rect 4723 22485 4753 22576
rect 4999 22485 5029 22576
rect 3065 22435 3105 22485
rect 3340 22435 3380 22485
rect 3615 22435 3655 22485
rect 3890 22435 3930 22485
rect 4165 22435 4205 22485
rect 4440 22435 4480 22485
rect 4715 22435 4755 22485
rect 4990 22435 5030 22485
rect 5275 22476 5305 22576
rect 5551 22476 5581 22576
rect 5827 22476 5857 22576
rect 6103 22476 6133 22576
rect 6379 22476 6409 22576
rect 6655 22476 6685 22576
rect 6931 22476 6961 22576
rect 7207 22476 7237 22576
rect 7483 22476 7513 22576
rect 7759 22476 7789 22576
rect 8035 22476 8065 22576
rect 8311 22476 8341 22576
rect 8587 22476 8617 22576
rect 8863 22476 8893 22576
rect 9139 22476 9169 22576
rect 9415 22476 9445 22576
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22476 11929 22576
rect 12175 22476 12205 22576
rect 12451 22476 12481 22576
rect 12727 22476 12757 22576
rect 13003 22476 13033 22576
rect 13279 22476 13309 22576
rect 13555 22476 13585 22576
rect 13831 22476 13861 22576
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 2710 22430 2760 22435
rect 2710 22390 2715 22430
rect 2755 22390 2760 22430
rect 2710 22385 2760 22390
rect 3060 22430 3110 22435
rect 3060 22390 3065 22430
rect 3105 22390 3110 22430
rect 3060 22385 3110 22390
rect 3335 22430 3385 22435
rect 3335 22390 3340 22430
rect 3380 22390 3385 22430
rect 3335 22385 3385 22390
rect 3610 22430 3660 22435
rect 3610 22390 3615 22430
rect 3655 22390 3660 22430
rect 3610 22385 3660 22390
rect 3885 22430 3935 22435
rect 3885 22390 3890 22430
rect 3930 22390 3935 22430
rect 3885 22385 3935 22390
rect 4160 22430 4210 22435
rect 4160 22390 4165 22430
rect 4205 22390 4210 22430
rect 4160 22385 4210 22390
rect 4435 22430 4485 22435
rect 4435 22390 4440 22430
rect 4480 22390 4485 22430
rect 4435 22385 4485 22390
rect 4710 22430 4760 22435
rect 4710 22390 4715 22430
rect 4755 22390 4760 22430
rect 4710 22385 4760 22390
rect 4985 22430 5035 22435
rect 4985 22390 4990 22430
rect 5030 22390 5035 22430
rect 4985 22385 5035 22390
rect 100 500 300 22076
rect 400 21980 600 22076
rect 2715 21985 2755 22385
rect 400 21940 405 21980
rect 445 21940 470 21980
rect 510 21940 535 21980
rect 575 21940 600 21980
rect 400 500 600 21940
rect 2710 21980 2760 21985
rect 2710 21940 2715 21980
rect 2755 21940 2760 21980
rect 2710 21935 2760 21940
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 19 nsew signal tristate
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 20 nsew signal tristate
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 21 nsew signal tristate
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 22 nsew signal tristate
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 23 nsew signal tristate
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 24 nsew signal tristate
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 25 nsew signal tristate
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 26 nsew signal tristate
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 27 nsew signal tristate
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 28 nsew signal tristate
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 29 nsew signal tristate
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 30 nsew signal tristate
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 31 nsew signal tristate
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 32 nsew signal tristate
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 33 nsew signal tristate
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 34 nsew signal tristate
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 35 nsew signal tristate
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 36 nsew signal tristate
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 37 nsew signal tristate
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 38 nsew signal tristate
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 39 nsew signal tristate
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 40 nsew signal tristate
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 41 nsew signal tristate
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 42 nsew signal tristate
flabel metal4 100 500 300 22076 1 FreeSans 1 0 0 0 VDPWR
port 43 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 1 0 0 0 VGND
port 44 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
