magic
tech sky130A
magscale 1 2
timestamp 1747494215
<< nwell >>
rect -40 260 9580 592
rect 455 -409 514 -88
rect 1104 -409 1129 -88
rect 1748 -409 1770 -88
rect 2388 -409 2413 -88
rect 2540 -100 2710 -78
rect 2540 -400 2630 -100
rect 2540 -420 2710 -400
rect 3234 -409 3270 -88
rect 3870 -409 3937 -88
rect 4543 -409 4568 -88
rect 5185 -406 5245 -88
rect 5394 -398 5460 -86
rect 5394 -406 5580 -398
rect 5185 -407 5580 -406
rect 6045 -407 6090 -86
rect 6700 -407 6754 -86
rect 7365 -407 7395 -86
rect 8013 -407 8068 -86
rect 8200 -90 8370 -80
rect 8200 -400 8300 -90
rect 5188 -410 5580 -407
rect 8200 -410 8370 -400
rect 8895 -407 8952 -86
rect 5400 -760 5570 -750
rect 540 -1081 630 -760
rect 1065 -1081 1182 -760
rect 1840 -1081 1940 -760
rect 2323 -1081 2417 -760
rect 2570 -1080 2630 -760
rect 2570 -1090 2750 -1080
rect 3337 -1081 3401 -760
rect 3838 -1081 3919 -760
rect 4634 -1081 4721 -760
rect 5156 -1081 5243 -760
rect 5400 -1080 5450 -760
rect 5400 -1090 5570 -1080
rect 6155 -1081 6239 -760
rect 6677 -1081 6752 -760
rect 7460 -1081 7541 -760
rect 7981 -1081 8064 -760
rect 8224 -1081 8276 -760
rect 8986 -1081 9131 -760
<< pwell >>
rect 1109 -49 1235 25
rect 1665 -48 1720 0
rect 1150 -650 1240 -450
rect 3810 -640 3990 -450
<< locali >>
rect 327 527 423 561
rect 1065 527 1217 561
rect 1619 527 1719 561
rect 2349 527 2453 561
rect 2532 527 2668 561
rect 3115 527 3233 561
rect 3866 527 3973 561
rect 4427 527 4530 561
rect 5170 527 5282 561
rect 5363 527 5481 561
rect 5928 527 6044 561
rect 6675 527 6792 561
rect 7246 527 7352 561
rect 7990 527 8104 561
rect 8184 527 8313 561
rect 8759 527 8894 561
rect -120 280 -40 300
rect -120 240 -100 280
rect -60 240 -40 280
rect -120 220 -40 240
rect 2030 249 2090 250
rect 2030 215 2047 249
rect 2081 215 2090 249
rect 2030 211 2090 215
rect 326 -17 424 17
rect 1061 -17 1221 17
rect 1618 -18 1720 17
rect 2348 -17 2457 17
rect 2526 -17 2661 17
rect 3115 -17 3235 17
rect 3863 -17 3973 17
rect 4417 -17 4534 17
rect 5170 -17 5285 17
rect 5359 -17 5483 17
rect 5925 -17 6047 17
rect 6678 -17 6794 17
rect 7237 -17 7354 17
rect 7981 -17 8104 17
rect 8178 -17 8315 17
rect 8768 -17 8894 17
rect 5110 -109 5280 -104
rect 1069 -143 1165 -109
rect 1712 -143 1842 -109
rect 2350 -143 2452 -109
rect 2523 -143 2664 -109
rect 3208 -143 3316 -109
rect 3828 -143 3974 -109
rect 4500 -143 4604 -109
rect 5110 -141 5282 -109
rect 5367 -141 5487 -107
rect 6027 -141 6121 -107
rect 6655 -141 6799 -107
rect 7337 -141 7433 -107
rect 7977 -141 8103 -107
rect 8183 -141 8314 -107
rect 8857 -141 8987 -107
rect 1712 -144 1759 -143
rect 5126 -653 5281 -651
rect 415 -687 524 -653
rect 1067 -687 1167 -653
rect 1711 -687 1843 -653
rect 2347 -687 2453 -653
rect 2533 -687 2665 -653
rect 3200 -687 3331 -653
rect 3830 -687 3976 -653
rect 4502 -687 4603 -653
rect 5126 -686 5285 -653
rect 5362 -685 5484 -651
rect 6027 -686 6126 -651
rect 6661 -685 6793 -651
rect 7333 -685 7433 -651
rect 7974 -685 8107 -651
rect 8189 -685 8313 -651
rect 8859 -685 8997 -651
rect 5126 -687 5281 -686
rect 2347 -688 2393 -687
rect 505 -815 670 -781
rect 1030 -815 1165 -781
rect 1804 -815 1925 -781
rect 2283 -815 2452 -781
rect 2537 -815 2660 -781
rect 3300 -815 3441 -781
rect 3803 -815 3973 -781
rect 4552 -815 4761 -781
rect 5124 -815 5283 -781
rect 5369 -815 5490 -781
rect 6119 -815 6276 -781
rect 6640 -815 6790 -781
rect 7431 -815 7580 -781
rect 7945 -815 8106 -781
rect 8187 -815 8318 -781
rect 8944 -815 9174 -781
rect 510 -1359 669 -1325
rect 1031 -1359 1165 -1325
rect 1803 -1359 1927 -1325
rect 2285 -1359 2452 -1325
rect 2528 -1359 2666 -1325
rect 3301 -1359 3439 -1325
rect 3804 -1359 3957 -1325
rect 4596 -1359 4762 -1325
rect 5124 -1359 5285 -1325
rect 5368 -1359 5484 -1325
rect 6120 -1359 6278 -1325
rect 6640 -1359 6789 -1325
rect 7431 -1359 7580 -1325
rect 7945 -1359 8101 -1325
rect 8186 -1359 8313 -1325
rect 8945 -1359 9174 -1325
<< viali >>
rect 8680 390 8720 430
rect -100 240 -60 280
rect 511 270 546 306
rect 1001 289 1035 323
rect 2295 289 2329 323
rect 3810 290 3850 330
rect 5095 307 5129 341
rect 6600 300 6640 340
rect 5880 260 5914 295
rect 7920 290 7960 330
rect 9460 290 9500 330
rect 80 220 120 260
rect 630 218 666 253
rect 1189 220 1223 255
rect 1375 215 1409 249
rect 1915 215 1950 251
rect 2047 215 2081 249
rect 2690 220 2730 260
rect 2873 223 2907 258
rect 3057 221 3092 255
rect 3320 215 3356 250
rect 3430 210 3470 250
rect 3990 220 4030 260
rect 4181 221 4215 255
rect 4370 200 4404 234
rect 4720 210 4760 250
rect 4865 218 4899 253
rect 5507 223 5541 258
rect 5690 220 5730 260
rect 6240 215 6274 249
rect 6375 215 6409 249
rect 6803 225 6840 260
rect 7001 221 7035 255
rect 7185 209 7219 245
rect 7433 215 7467 249
rect 7550 217 7584 252
rect 8339 221 8373 255
rect 8525 215 8559 249
rect 9092 215 9126 249
rect 9220 210 9260 250
rect 267 153 301 187
rect 1560 140 1600 180
rect -113 -256 -79 -220
rect 3974 -260 4014 -220
rect 8334 -290 8370 -251
rect 5500 -390 5540 -350
rect 83 -457 128 -417
rect 348 -455 382 -421
rect 1388 -455 1422 -421
rect 1505 -455 1540 -421
rect 1644 -455 1678 -421
rect 2882 -453 2916 -419
rect 3138 -455 3172 -421
rect 4192 -455 4226 -421
rect 4438 -455 4472 -421
rect 5690 -450 5730 -408
rect 5820 -460 5860 -420
rect 5958 -453 5992 -419
rect 7020 -450 7060 -410
rect 7140 -450 7180 -410
rect 7268 -453 7302 -419
rect 8540 -450 8580 -410
rect 8790 -453 8824 -419
rect 260 -570 300 -530
rect 1199 -575 1233 -541
rect 2680 -560 2720 -520
rect 3055 -580 3090 -543
rect 4350 -570 4390 -530
rect 6810 -570 6850 -530
rect 8706 -567 8741 -533
rect 440 -970 480 -930
rect 1731 -967 1765 -933
rect 3239 -1053 3273 -1019
rect 4540 -1060 4580 -1020
rect 6050 -1050 6090 -1010
rect 8400 -1070 8435 -1036
rect 8890 -1050 8930 -1010
rect -45 -1127 -11 -1093
rect 70 -1127 104 -1093
rect 1250 -1140 1290 -1090
rect 1364 -1127 1398 -1093
rect 2747 -1130 2783 -1093
rect 2860 -1127 2894 -1093
rect 4053 -1127 4087 -1093
rect 4170 -1127 4204 -1093
rect 5563 -1127 5597 -1093
rect 5680 -1127 5714 -1093
rect 6873 -1127 6907 -1093
rect 6990 -1127 7024 -1093
rect 8510 -1127 8544 -1093
rect 7289 -1230 7323 -1193
<< metal1 >>
rect 325 496 426 592
rect 1063 496 1218 592
rect 1615 496 1720 592
rect 2354 496 2456 592
rect 2537 496 2661 592
rect 3110 496 3238 592
rect 3851 496 3977 592
rect 4423 496 4532 592
rect 5167 496 5282 592
rect 5367 496 5484 592
rect 5934 496 6044 592
rect 6679 496 6791 592
rect 7240 496 7354 592
rect 7987 496 8105 592
rect 8188 496 8312 592
rect 8765 496 8898 592
rect 8650 450 8740 460
rect 8650 380 8660 450
rect 8730 380 8740 450
rect 8650 370 8740 380
rect 5070 350 5150 360
rect 2270 340 2350 350
rect 980 330 1060 340
rect 470 320 559 330
rect -120 290 -40 300
rect -120 230 -110 290
rect -50 230 -40 290
rect -120 220 -40 230
rect 60 272 140 290
rect 60 210 70 272
rect 130 210 140 272
rect 470 260 480 320
rect 540 306 559 320
rect 546 270 559 306
rect 610 280 690 290
rect 610 270 620 280
rect 540 260 559 270
rect 470 250 550 260
rect 600 220 620 270
rect 680 220 690 280
rect 980 270 990 330
rect 1050 270 1060 330
rect 2270 280 2280 340
rect 2340 280 2350 340
rect 3780 340 3860 350
rect 3780 280 3790 340
rect 3850 280 3860 340
rect 5070 290 5080 350
rect 5140 290 5150 350
rect 6580 350 6660 360
rect 5860 310 5940 320
rect 5070 280 5150 290
rect 5490 280 5570 290
rect 1900 270 1980 280
rect 2270 270 2350 280
rect 2680 270 2760 280
rect 980 260 1060 270
rect 1150 260 1230 270
rect 600 218 630 220
rect 666 218 690 220
rect 600 210 690 218
rect 1150 200 1160 260
rect 1220 255 1230 260
rect 1223 220 1230 255
rect 1220 200 1230 220
rect 230 190 320 200
rect 1150 190 1230 200
rect 1350 260 1430 270
rect 1350 200 1360 260
rect 1420 200 1430 260
rect 1900 210 1910 270
rect 1970 210 1980 270
rect 1900 200 1980 210
rect 2020 260 2100 270
rect 2020 200 2030 260
rect 2090 200 2100 260
rect 2680 210 2690 270
rect 2750 210 2760 270
rect 2680 200 2760 210
rect 2850 270 2930 280
rect 3410 270 3490 280
rect 3780 270 3860 280
rect 3960 270 4040 280
rect 2850 210 2860 270
rect 2920 210 2930 270
rect 1350 190 1430 200
rect 1540 190 1620 200
rect 2020 190 2100 200
rect 2850 190 2930 210
rect 3050 260 3130 270
rect 3313 260 3362 270
rect 3050 255 3060 260
rect 3050 221 3057 255
rect 3050 200 3060 221
rect 3120 200 3130 260
rect 3050 190 3130 200
rect 3280 250 3362 260
rect 3280 190 3290 250
rect 3356 215 3362 250
rect 3350 199 3362 215
rect 3410 210 3420 270
rect 3480 210 3490 270
rect 3410 200 3490 210
rect 3960 210 3970 270
rect 4030 210 4040 270
rect 4167 260 4235 265
rect 3960 200 4040 210
rect 4160 255 4240 260
rect 4160 250 4181 255
rect 4215 250 4240 255
rect 3350 190 3360 199
rect 4160 190 4170 250
rect 4230 190 4240 250
rect 230 130 250 190
rect 310 130 320 190
rect 230 120 320 130
rect 1540 130 1550 190
rect 1610 130 1620 190
rect 4160 180 4240 190
rect 4360 250 4440 260
rect 4360 190 4370 250
rect 4430 190 4440 250
rect 4700 210 4720 270
rect 4780 210 4800 270
rect 4700 200 4800 210
rect 4840 260 4920 271
rect 4360 180 4440 190
rect 4840 199 4850 260
rect 4910 199 4920 260
rect 5490 220 5500 280
rect 5560 220 5570 280
rect 5490 210 5570 220
rect 5670 270 5760 280
rect 5670 210 5680 270
rect 5740 210 5760 270
rect 5860 250 5870 310
rect 5930 250 5940 310
rect 6580 290 6590 350
rect 6650 290 6660 350
rect 9440 340 9520 350
rect 6580 280 6660 290
rect 7900 330 7980 340
rect 7520 270 7600 280
rect 6780 260 6860 270
rect 5860 240 5940 250
rect 6200 250 6330 260
rect 4840 179 4920 199
rect 5670 170 5760 210
rect 6200 190 6220 250
rect 6280 190 6330 250
rect 6200 170 6330 190
rect 6360 250 6440 260
rect 6360 190 6370 250
rect 6430 190 6440 250
rect 6780 200 6790 260
rect 6850 200 6860 260
rect 6780 190 6860 200
rect 6980 260 7060 270
rect 7520 260 7530 270
rect 6980 200 6990 260
rect 7050 200 7060 260
rect 6980 190 7060 200
rect 7170 250 7250 260
rect 7170 190 7180 250
rect 7240 190 7250 250
rect 6360 180 6440 190
rect 7170 180 7250 190
rect 7399 250 7480 260
rect 7399 190 7410 250
rect 7470 190 7480 250
rect 7510 210 7530 260
rect 7590 260 7600 270
rect 7900 270 7910 330
rect 7970 270 7980 330
rect 7900 260 7980 270
rect 8290 290 8380 310
rect 7590 210 7630 260
rect 8290 230 8300 290
rect 8360 270 8380 290
rect 9440 280 9450 340
rect 9510 280 9520 340
rect 8360 255 8399 270
rect 8290 221 8339 230
rect 8373 221 8399 255
rect 8290 210 8399 221
rect 8500 260 8590 270
rect 7520 200 7600 210
rect 8500 200 8510 260
rect 8570 200 8590 260
rect 8500 190 8590 200
rect 9050 260 9180 270
rect 9050 200 9060 260
rect 9120 249 9180 260
rect 9126 215 9180 249
rect 9120 200 9180 215
rect 9050 190 9180 200
rect 9210 260 9310 280
rect 9440 270 9520 280
rect 9210 200 9220 260
rect 9280 200 9310 260
rect 9210 190 9310 200
rect 7399 170 7480 190
rect 1540 120 1620 130
rect 317 -48 320 48
rect 323 -48 427 48
rect 1063 -49 1223 48
rect 1615 -48 1720 48
rect 2352 17 2461 48
rect 2348 -17 2461 17
rect 2352 -49 2461 -17
rect 2535 -48 2666 48
rect 3111 -48 3238 48
rect 3867 -48 3973 48
rect 4423 -14 4532 48
rect 4422 -48 4534 -14
rect 5166 -48 5285 48
rect 5365 -48 5486 48
rect 5933 -48 6045 48
rect 6675 -48 6794 48
rect 7244 -48 7357 48
rect 7986 -48 8108 48
rect 8185 -48 8314 48
rect 8761 -48 8894 48
rect 417 -174 521 -78
rect 1066 -174 1167 -78
rect 1708 -174 1846 -78
rect 2345 -174 2454 -78
rect 2532 -174 2664 -78
rect 3200 -174 3310 -78
rect 3835 -174 3976 -78
rect 4504 -174 4606 -78
rect 5110 -172 5283 -78
rect 5361 -172 5487 -76
rect 6023 -172 6124 -76
rect 6665 -172 6794 -76
rect 7334 -172 7431 -76
rect 7974 -172 8104 -76
rect 8186 -172 8313 -76
rect 8845 -172 8988 -76
rect -130 -220 -50 -210
rect -130 -280 -120 -220
rect -60 -280 -50 -220
rect -130 -290 -50 -280
rect 3960 -220 4040 -210
rect 3960 -280 3970 -220
rect 4030 -280 4040 -220
rect 3960 -290 4040 -280
rect 8310 -230 8390 -220
rect 8310 -290 8320 -230
rect 8380 -290 8390 -230
rect 8310 -300 8390 -290
rect 5480 -340 5560 -330
rect 50 -400 130 -390
rect 340 -400 420 -390
rect 50 -460 60 -400
rect 120 -417 140 -400
rect 128 -457 140 -417
rect 120 -460 140 -457
rect 50 -470 140 -460
rect 340 -421 350 -400
rect 340 -455 348 -421
rect 340 -460 350 -455
rect 410 -460 420 -400
rect 340 -470 420 -460
rect 1370 -400 1450 -390
rect 1370 -460 1380 -400
rect 1440 -460 1450 -400
rect 1370 -470 1450 -460
rect 1490 -400 1570 -380
rect 2850 -390 2930 -380
rect 1490 -460 1500 -400
rect 1560 -460 1570 -400
rect 1490 -470 1570 -460
rect 1630 -400 1710 -390
rect 1630 -460 1640 -400
rect 1700 -460 1710 -400
rect 2850 -450 2860 -390
rect 2920 -450 2930 -390
rect 2850 -453 2882 -450
rect 2916 -453 2930 -450
rect 2850 -460 2930 -453
rect 3130 -400 3210 -390
rect 3130 -421 3140 -400
rect 3130 -455 3138 -421
rect 3130 -460 3140 -455
rect 3200 -460 3210 -400
rect 1630 -470 1710 -460
rect 3130 -470 3210 -460
rect 4170 -400 4250 -390
rect 4170 -460 4180 -400
rect 4240 -460 4250 -400
rect 4170 -470 4250 -460
rect 4430 -400 4510 -390
rect 4430 -421 4440 -400
rect 4430 -455 4438 -421
rect 4430 -460 4440 -455
rect 4500 -460 4510 -400
rect 5480 -400 5490 -340
rect 5550 -400 5560 -340
rect 5480 -410 5560 -400
rect 5670 -390 5750 -380
rect 5670 -450 5680 -390
rect 5740 -450 5750 -390
rect 5670 -460 5750 -450
rect 5800 -400 5880 -390
rect 5800 -460 5810 -400
rect 5870 -460 5880 -400
rect 4430 -470 4510 -460
rect 5800 -470 5880 -460
rect 5940 -399 6020 -390
rect 5940 -460 5950 -399
rect 6010 -460 6020 -399
rect 5940 -470 6020 -460
rect 6990 -400 7070 -390
rect 6990 -460 7000 -400
rect 7060 -460 7070 -400
rect 6990 -470 7070 -460
rect 7120 -400 7200 -390
rect 7120 -460 7130 -400
rect 7190 -460 7200 -400
rect 7120 -470 7200 -460
rect 7260 -400 7340 -390
rect 7260 -419 7270 -400
rect 7260 -453 7268 -419
rect 7260 -460 7270 -453
rect 7330 -460 7340 -400
rect 7260 -470 7340 -460
rect 8520 -400 8600 -390
rect 8520 -460 8530 -400
rect 8590 -460 8600 -400
rect 8520 -470 8600 -460
rect 8780 -410 8860 -400
rect 8780 -470 8790 -410
rect 8850 -470 8860 -410
rect 8780 -480 8860 -470
rect 2650 -510 2730 -500
rect 8670 -510 8750 -500
rect 250 -520 340 -510
rect 250 -580 260 -520
rect 320 -580 340 -520
rect 250 -590 340 -580
rect 1160 -520 1240 -510
rect 1160 -580 1170 -520
rect 1230 -541 1240 -520
rect 1233 -575 1240 -541
rect 1230 -580 1240 -575
rect 2650 -570 2660 -510
rect 2720 -570 2730 -510
rect 2650 -580 2730 -570
rect 3030 -520 3110 -510
rect 3030 -580 3040 -520
rect 3100 -580 3110 -520
rect 1160 -590 1240 -580
rect 3030 -590 3110 -580
rect 4320 -520 4400 -510
rect 4320 -580 4330 -520
rect 4390 -580 4400 -520
rect 4320 -590 4400 -580
rect 6780 -520 6860 -510
rect 6780 -580 6790 -520
rect 6850 -580 6860 -520
rect 8670 -570 8680 -510
rect 8740 -533 8750 -510
rect 8741 -567 8750 -533
rect 8740 -570 8750 -567
rect 8670 -580 8750 -570
rect 6780 -590 6860 -580
rect 417 -718 523 -622
rect 1065 -718 1168 -622
rect 1709 -718 1843 -622
rect 2352 -718 2453 -622
rect 2535 -718 2666 -622
rect 3204 -718 3326 -622
rect 3834 -718 3976 -622
rect 4484 -718 4604 -622
rect 5144 -720 5283 -620
rect 5365 -716 5487 -620
rect 6024 -716 6125 -620
rect 6666 -716 6795 -620
rect 7336 -716 7436 -620
rect 7977 -716 8107 -620
rect 8186 -716 8315 -620
rect 8856 -716 8992 -620
rect 508 -846 670 -750
rect 1028 -846 1166 -750
rect 1803 -846 1925 -750
rect 2288 -846 2452 -750
rect 2535 -846 2662 -750
rect 3297 -846 3443 -750
rect 3800 -846 3974 -750
rect 4574 -846 4766 -750
rect 5120 -846 5284 -750
rect 5366 -846 5484 -750
rect 6115 -846 6278 -750
rect 6637 -846 6791 -750
rect 7429 -846 7581 -750
rect 7943 -770 8112 -750
rect 7943 -840 8110 -770
rect 7943 -846 8112 -840
rect 8181 -846 8314 -750
rect 8937 -846 9175 -750
rect 430 -920 510 -910
rect 430 -980 440 -920
rect 500 -980 510 -920
rect 430 -990 510 -980
rect 1720 -920 1800 -910
rect 1720 -980 1729 -920
rect 1789 -980 1800 -920
rect 1720 -990 1800 -980
rect 6030 -970 6050 -910
rect 6110 -970 6120 -910
rect 3220 -1000 3300 -990
rect 3220 -1060 3230 -1000
rect 3290 -1060 3300 -1000
rect 4520 -1000 4600 -990
rect 4520 -1060 4530 -1000
rect 4590 -1060 4600 -1000
rect 6030 -1010 6120 -970
rect 8870 -1000 8950 -990
rect 6030 -1050 6050 -1010
rect 6090 -1050 6120 -1010
rect 2840 -1070 2920 -1060
rect 3220 -1070 3300 -1060
rect 4020 -1070 4100 -1060
rect -70 -1080 10 -1070
rect -70 -1140 -60 -1080
rect 0 -1140 10 -1080
rect -70 -1150 10 -1140
rect 50 -1080 130 -1070
rect 1340 -1080 1420 -1070
rect 50 -1141 60 -1080
rect 120 -1141 130 -1080
rect 50 -1150 130 -1141
rect 1230 -1088 1310 -1080
rect 1230 -1150 1240 -1088
rect 1300 -1150 1310 -1088
rect 1340 -1140 1350 -1080
rect 1410 -1140 1420 -1080
rect 1340 -1150 1420 -1140
rect 2720 -1080 2800 -1070
rect 2720 -1140 2730 -1080
rect 2790 -1140 2800 -1080
rect 2840 -1130 2850 -1070
rect 2910 -1130 2920 -1070
rect 2840 -1140 2920 -1130
rect 4020 -1130 4030 -1070
rect 4090 -1130 4100 -1070
rect 4020 -1140 4100 -1130
rect 4150 -1070 4230 -1060
rect 4520 -1070 4600 -1060
rect 5670 -1070 5750 -1060
rect 6030 -1070 6120 -1050
rect 8370 -1010 8450 -1000
rect 8370 -1070 8380 -1010
rect 8440 -1070 8450 -1010
rect 8870 -1060 8880 -1000
rect 8940 -1060 8950 -1000
rect 4150 -1130 4160 -1070
rect 4220 -1130 4230 -1070
rect 4150 -1140 4230 -1130
rect 5540 -1080 5620 -1070
rect 5540 -1140 5550 -1080
rect 5610 -1140 5620 -1080
rect 5670 -1130 5680 -1070
rect 5740 -1130 5750 -1070
rect 5670 -1140 5750 -1130
rect 6850 -1080 6930 -1070
rect 6850 -1140 6860 -1080
rect 6920 -1140 6930 -1080
rect 2720 -1150 2800 -1140
rect 5540 -1150 5620 -1140
rect 6850 -1150 6930 -1140
rect 6970 -1080 7050 -1070
rect 8370 -1080 8450 -1070
rect 8490 -1070 8570 -1060
rect 8870 -1070 8950 -1060
rect 6970 -1140 6980 -1080
rect 7040 -1140 7050 -1080
rect 8490 -1130 8500 -1070
rect 8560 -1130 8570 -1070
rect 8490 -1140 8570 -1130
rect 6970 -1150 7050 -1140
rect 1230 -1160 1310 -1150
rect 7270 -1170 7360 -1160
rect 7270 -1193 7290 -1170
rect 7270 -1230 7289 -1193
rect 7350 -1230 7360 -1170
rect 7270 -1240 7360 -1230
rect 7270 -1250 7309 -1240
rect 507 -1390 670 -1294
rect 1025 -1390 1168 -1294
rect 1801 -1390 1929 -1294
rect 2288 -1390 2452 -1294
rect 2534 -1390 2665 -1294
rect 3298 -1390 3442 -1294
rect 3802 -1390 3957 -1294
rect 4594 -1390 4760 -1294
rect 5121 -1300 5292 -1294
rect 5121 -1370 5290 -1300
rect 5121 -1390 5292 -1370
rect 5364 -1390 5488 -1294
rect 6118 -1390 6276 -1294
rect 6636 -1390 6791 -1294
rect 7430 -1390 7579 -1294
rect 7944 -1390 8101 -1294
rect 8188 -1390 8316 -1294
rect 8944 -1390 9170 -1294
<< via1 >>
rect 8110 510 8180 580
rect 8660 430 8730 450
rect 8660 390 8680 430
rect 8680 390 8720 430
rect 8720 390 8730 430
rect 8660 380 8730 390
rect -110 280 -50 290
rect -110 240 -100 280
rect -100 240 -60 280
rect -60 240 -50 280
rect -110 230 -50 240
rect 70 260 130 272
rect 70 220 80 260
rect 80 220 120 260
rect 120 220 130 260
rect 70 210 130 220
rect 480 306 540 320
rect 480 270 511 306
rect 511 270 540 306
rect 480 260 540 270
rect 620 253 680 280
rect 620 220 630 253
rect 630 220 666 253
rect 666 220 680 253
rect 990 323 1050 330
rect 990 289 1001 323
rect 1001 289 1035 323
rect 1035 289 1050 323
rect 990 270 1050 289
rect 2280 323 2340 340
rect 2280 289 2295 323
rect 2295 289 2329 323
rect 2329 289 2340 323
rect 2280 280 2340 289
rect 3790 330 3850 340
rect 3790 290 3810 330
rect 3810 290 3850 330
rect 3790 280 3850 290
rect 5080 341 5140 350
rect 5080 307 5095 341
rect 5095 307 5129 341
rect 5129 307 5140 341
rect 5080 290 5140 307
rect 1160 255 1220 260
rect 1160 220 1189 255
rect 1189 220 1220 255
rect 1160 200 1220 220
rect 1360 249 1420 260
rect 1360 215 1375 249
rect 1375 215 1409 249
rect 1409 215 1420 249
rect 1360 200 1420 215
rect 1910 251 1970 270
rect 1910 215 1915 251
rect 1915 215 1950 251
rect 1950 215 1970 251
rect 1910 210 1970 215
rect 2030 249 2090 260
rect 2030 215 2047 249
rect 2047 215 2081 249
rect 2081 215 2090 249
rect 2030 200 2090 215
rect 2690 260 2750 270
rect 2690 220 2730 260
rect 2730 220 2750 260
rect 2690 210 2750 220
rect 2860 258 2920 270
rect 2860 223 2873 258
rect 2873 223 2907 258
rect 2907 223 2920 258
rect 2860 210 2920 223
rect 3060 255 3120 260
rect 3060 221 3092 255
rect 3092 221 3120 255
rect 3060 200 3120 221
rect 3290 215 3320 250
rect 3320 215 3350 250
rect 3290 190 3350 215
rect 3420 250 3480 270
rect 3420 210 3430 250
rect 3430 210 3470 250
rect 3470 210 3480 250
rect 3970 260 4030 270
rect 3970 220 3990 260
rect 3990 220 4030 260
rect 3970 210 4030 220
rect 4170 221 4181 250
rect 4181 221 4215 250
rect 4215 221 4230 250
rect 4170 190 4230 221
rect 250 187 310 190
rect 250 153 267 187
rect 267 153 301 187
rect 301 153 310 187
rect 250 130 310 153
rect 1550 180 1610 190
rect 1550 140 1560 180
rect 1560 140 1600 180
rect 1600 140 1610 180
rect 1550 130 1610 140
rect 4370 234 4430 250
rect 4370 200 4404 234
rect 4404 200 4430 234
rect 4370 190 4430 200
rect 4720 250 4780 270
rect 4720 210 4760 250
rect 4760 210 4780 250
rect 4850 253 4910 260
rect 4850 218 4865 253
rect 4865 218 4899 253
rect 4899 218 4910 253
rect 4850 199 4910 218
rect 5500 258 5560 280
rect 5500 223 5507 258
rect 5507 223 5541 258
rect 5541 223 5560 258
rect 5500 220 5560 223
rect 5680 260 5740 270
rect 5680 220 5690 260
rect 5690 220 5730 260
rect 5730 220 5740 260
rect 5680 210 5740 220
rect 5870 295 5930 310
rect 5870 260 5880 295
rect 5880 260 5914 295
rect 5914 260 5930 295
rect 5870 250 5930 260
rect 6590 340 6650 350
rect 6590 300 6600 340
rect 6600 300 6640 340
rect 6640 300 6650 340
rect 6590 290 6650 300
rect 6220 249 6280 250
rect 6220 215 6240 249
rect 6240 215 6274 249
rect 6274 215 6280 249
rect 6220 190 6280 215
rect 6370 249 6430 250
rect 6370 215 6375 249
rect 6375 215 6409 249
rect 6409 215 6430 249
rect 6370 190 6430 215
rect 6790 225 6803 260
rect 6803 225 6840 260
rect 6840 225 6850 260
rect 6790 200 6850 225
rect 6990 255 7050 260
rect 6990 221 7001 255
rect 7001 221 7035 255
rect 7035 221 7050 255
rect 6990 200 7050 221
rect 7180 245 7240 250
rect 7180 209 7185 245
rect 7185 209 7219 245
rect 7219 209 7240 245
rect 7180 190 7240 209
rect 7410 249 7470 250
rect 7410 215 7433 249
rect 7433 215 7467 249
rect 7467 215 7470 249
rect 7410 190 7470 215
rect 7530 252 7590 270
rect 7910 290 7920 330
rect 7920 290 7960 330
rect 7960 290 7970 330
rect 7910 270 7970 290
rect 7530 217 7550 252
rect 7550 217 7584 252
rect 7584 217 7590 252
rect 7530 210 7590 217
rect 8300 255 8360 290
rect 9450 330 9510 340
rect 9450 290 9460 330
rect 9460 290 9500 330
rect 9500 290 9510 330
rect 9450 280 9510 290
rect 8300 230 8339 255
rect 8339 230 8360 255
rect 8510 249 8570 260
rect 8510 215 8525 249
rect 8525 215 8559 249
rect 8559 215 8570 249
rect 8510 200 8570 215
rect 9060 249 9120 260
rect 9060 215 9092 249
rect 9092 215 9120 249
rect 9060 200 9120 215
rect 9220 250 9280 260
rect 9220 210 9260 250
rect 9260 210 9280 250
rect 9220 200 9280 210
rect 5290 -30 5360 40
rect 8110 -170 8180 -100
rect -120 -256 -113 -220
rect -113 -256 -79 -220
rect -79 -256 -60 -220
rect -120 -280 -60 -256
rect 3970 -260 3974 -220
rect 3974 -260 4014 -220
rect 4014 -260 4030 -220
rect 3970 -280 4030 -260
rect 8320 -251 8380 -230
rect 8320 -290 8334 -251
rect 8334 -290 8370 -251
rect 8370 -290 8380 -251
rect 60 -417 120 -400
rect 60 -457 83 -417
rect 83 -457 120 -417
rect 60 -460 120 -457
rect 350 -421 410 -400
rect 350 -455 382 -421
rect 382 -455 410 -421
rect 350 -460 410 -455
rect 1380 -421 1440 -400
rect 1380 -455 1388 -421
rect 1388 -455 1422 -421
rect 1422 -455 1440 -421
rect 1380 -460 1440 -455
rect 1500 -421 1560 -400
rect 1500 -455 1505 -421
rect 1505 -455 1540 -421
rect 1540 -455 1560 -421
rect 1500 -460 1560 -455
rect 1640 -421 1700 -400
rect 1640 -455 1644 -421
rect 1644 -455 1678 -421
rect 1678 -455 1700 -421
rect 1640 -460 1700 -455
rect 2860 -419 2920 -390
rect 2860 -450 2882 -419
rect 2882 -450 2916 -419
rect 2916 -450 2920 -419
rect 3140 -421 3200 -400
rect 3140 -455 3172 -421
rect 3172 -455 3200 -421
rect 3140 -460 3200 -455
rect 4180 -421 4240 -400
rect 4180 -455 4192 -421
rect 4192 -455 4226 -421
rect 4226 -455 4240 -421
rect 4180 -460 4240 -455
rect 4440 -421 4500 -400
rect 4440 -455 4472 -421
rect 4472 -455 4500 -421
rect 4440 -460 4500 -455
rect 5490 -350 5550 -340
rect 5490 -390 5500 -350
rect 5500 -390 5540 -350
rect 5540 -390 5550 -350
rect 5490 -400 5550 -390
rect 5680 -408 5740 -390
rect 5680 -450 5690 -408
rect 5690 -450 5730 -408
rect 5730 -450 5740 -408
rect 5810 -420 5870 -400
rect 5810 -460 5820 -420
rect 5820 -460 5860 -420
rect 5860 -460 5870 -420
rect 5950 -419 6010 -399
rect 5950 -453 5958 -419
rect 5958 -453 5992 -419
rect 5992 -453 6010 -419
rect 5950 -460 6010 -453
rect 7000 -410 7060 -400
rect 7000 -450 7020 -410
rect 7020 -450 7060 -410
rect 7000 -460 7060 -450
rect 7130 -410 7190 -400
rect 7130 -450 7140 -410
rect 7140 -450 7180 -410
rect 7180 -450 7190 -410
rect 7130 -460 7190 -450
rect 7270 -419 7330 -400
rect 7270 -453 7302 -419
rect 7302 -453 7330 -419
rect 7270 -460 7330 -453
rect 8530 -410 8590 -400
rect 8530 -450 8540 -410
rect 8540 -450 8580 -410
rect 8580 -450 8590 -410
rect 8530 -460 8590 -450
rect 8790 -419 8850 -410
rect 8790 -453 8824 -419
rect 8824 -453 8850 -419
rect 8790 -470 8850 -453
rect 260 -530 320 -520
rect 260 -570 300 -530
rect 300 -570 320 -530
rect 260 -580 320 -570
rect 1170 -541 1230 -520
rect 1170 -575 1199 -541
rect 1199 -575 1230 -541
rect 1170 -580 1230 -575
rect 2660 -520 2720 -510
rect 2660 -560 2680 -520
rect 2680 -560 2720 -520
rect 2660 -570 2720 -560
rect 3040 -543 3100 -520
rect 3040 -580 3055 -543
rect 3055 -580 3090 -543
rect 3090 -580 3100 -543
rect 4330 -530 4390 -520
rect 4330 -570 4350 -530
rect 4350 -570 4390 -530
rect 4330 -580 4390 -570
rect 6790 -530 6850 -520
rect 6790 -570 6810 -530
rect 6810 -570 6850 -530
rect 6790 -580 6850 -570
rect 8680 -533 8740 -510
rect 8680 -567 8706 -533
rect 8706 -567 8740 -533
rect 8680 -570 8740 -567
rect 5290 -700 5360 -630
rect 8110 -840 8180 -770
rect 440 -930 500 -920
rect 440 -970 480 -930
rect 480 -970 500 -930
rect 440 -980 500 -970
rect 1729 -933 1789 -920
rect 1729 -967 1731 -933
rect 1731 -967 1765 -933
rect 1765 -967 1789 -933
rect 1729 -980 1789 -967
rect 6050 -970 6110 -910
rect 3230 -1019 3290 -1000
rect 3230 -1053 3239 -1019
rect 3239 -1053 3273 -1019
rect 3273 -1053 3290 -1019
rect 3230 -1060 3290 -1053
rect 4530 -1020 4590 -1000
rect 4530 -1060 4540 -1020
rect 4540 -1060 4580 -1020
rect 4580 -1060 4590 -1020
rect -60 -1093 0 -1080
rect -60 -1127 -45 -1093
rect -45 -1127 -11 -1093
rect -11 -1127 0 -1093
rect -60 -1140 0 -1127
rect 60 -1093 120 -1080
rect 60 -1127 70 -1093
rect 70 -1127 104 -1093
rect 104 -1127 120 -1093
rect 60 -1141 120 -1127
rect 1240 -1090 1300 -1088
rect 1240 -1140 1250 -1090
rect 1250 -1140 1290 -1090
rect 1290 -1140 1300 -1090
rect 1240 -1150 1300 -1140
rect 1350 -1093 1410 -1080
rect 1350 -1127 1364 -1093
rect 1364 -1127 1398 -1093
rect 1398 -1127 1410 -1093
rect 1350 -1140 1410 -1127
rect 2730 -1093 2790 -1080
rect 2730 -1130 2747 -1093
rect 2747 -1130 2783 -1093
rect 2783 -1130 2790 -1093
rect 2730 -1140 2790 -1130
rect 2850 -1093 2910 -1070
rect 2850 -1127 2860 -1093
rect 2860 -1127 2894 -1093
rect 2894 -1127 2910 -1093
rect 2850 -1130 2910 -1127
rect 4030 -1093 4090 -1070
rect 4030 -1127 4053 -1093
rect 4053 -1127 4087 -1093
rect 4087 -1127 4090 -1093
rect 4030 -1130 4090 -1127
rect 8380 -1036 8440 -1010
rect 8380 -1070 8400 -1036
rect 8400 -1070 8435 -1036
rect 8435 -1070 8440 -1036
rect 8880 -1010 8940 -1000
rect 8880 -1050 8890 -1010
rect 8890 -1050 8930 -1010
rect 8930 -1050 8940 -1010
rect 8880 -1060 8940 -1050
rect 4160 -1093 4220 -1070
rect 4160 -1127 4170 -1093
rect 4170 -1127 4204 -1093
rect 4204 -1127 4220 -1093
rect 4160 -1130 4220 -1127
rect 5550 -1093 5610 -1080
rect 5550 -1127 5563 -1093
rect 5563 -1127 5597 -1093
rect 5597 -1127 5610 -1093
rect 5550 -1140 5610 -1127
rect 5680 -1093 5740 -1070
rect 5680 -1127 5714 -1093
rect 5714 -1127 5740 -1093
rect 5680 -1130 5740 -1127
rect 6860 -1093 6920 -1080
rect 6860 -1127 6873 -1093
rect 6873 -1127 6907 -1093
rect 6907 -1127 6920 -1093
rect 6860 -1140 6920 -1127
rect 6980 -1093 7040 -1080
rect 6980 -1127 6990 -1093
rect 6990 -1127 7024 -1093
rect 7024 -1127 7040 -1093
rect 6980 -1140 7040 -1127
rect 8500 -1093 8560 -1070
rect 8500 -1127 8510 -1093
rect 8510 -1127 8544 -1093
rect 8544 -1127 8560 -1093
rect 8500 -1130 8560 -1127
rect 7290 -1193 7350 -1170
rect 7290 -1230 7323 -1193
rect 7323 -1230 7350 -1193
rect 5290 -1370 5360 -1300
<< metal2 >>
rect 8100 580 8190 590
rect 2680 500 2760 530
rect -130 440 -30 460
rect -130 380 -110 440
rect -50 380 -30 440
rect -130 360 -30 380
rect 610 440 690 460
rect 670 380 690 440
rect -120 290 -40 360
rect 470 320 570 330
rect -120 230 -110 290
rect -50 230 -40 290
rect -120 220 -40 230
rect 60 272 140 290
rect 60 210 70 272
rect 130 210 140 272
rect 470 260 480 320
rect 540 260 570 320
rect 470 250 570 260
rect 70 180 150 210
rect 60 160 150 180
rect 60 100 70 160
rect 130 100 150 160
rect 230 190 320 200
rect 230 130 250 190
rect 310 130 320 190
rect 490 180 570 250
rect 610 280 690 380
rect 1140 440 1230 460
rect 1140 380 1160 440
rect 1220 380 1230 440
rect 1140 360 1230 380
rect 610 220 620 280
rect 680 220 690 280
rect 980 330 1060 340
rect 980 270 990 330
rect 980 260 1060 270
rect 1150 260 1230 360
rect 1900 430 1990 460
rect 1900 370 1910 430
rect 1970 370 1990 430
rect 1900 290 1990 370
rect 2680 440 2690 500
rect 2750 440 2760 500
rect 1890 270 1990 290
rect 2270 340 2350 350
rect 2270 280 2280 340
rect 2340 280 2350 340
rect 2270 270 2350 280
rect 2680 270 2760 440
rect 3410 500 3490 530
rect 3410 440 3420 500
rect 3480 440 3490 500
rect 8100 510 8110 580
rect 8180 510 8190 580
rect 5490 460 5570 480
rect 610 210 690 220
rect 1150 200 1160 260
rect 1220 200 1230 260
rect 1150 190 1230 200
rect 1350 260 1430 270
rect 1350 200 1360 260
rect 1420 200 1430 260
rect 1890 210 1910 270
rect 1970 210 1990 270
rect 230 120 320 130
rect 480 160 570 180
rect 1350 170 1430 200
rect 1540 190 1620 200
rect 1890 190 1990 210
rect 2020 260 2100 270
rect 2020 200 2030 260
rect 2090 200 2100 260
rect 2680 210 2690 270
rect 2750 210 2760 270
rect 2680 200 2760 210
rect 2850 270 2930 279
rect 2850 210 2860 270
rect 2920 210 2930 270
rect 60 80 150 100
rect 250 20 310 120
rect 480 100 500 160
rect 560 100 570 160
rect 480 80 570 100
rect 1340 150 1440 170
rect 1340 90 1360 150
rect 1420 90 1440 150
rect 1340 70 1440 90
rect 1540 130 1550 190
rect 1610 130 1620 190
rect 50 10 130 20
rect 50 -50 60 10
rect 120 -50 130 10
rect 50 -60 130 -50
rect 230 10 310 20
rect 230 -50 240 10
rect 300 -50 310 10
rect 230 -60 310 -50
rect 1370 -60 1450 -50
rect -130 -220 -50 -210
rect -130 -280 -120 -220
rect -60 -280 -50 -220
rect -130 -290 -50 -280
rect 50 -370 110 -60
rect 1370 -120 1380 -60
rect 1440 -120 1450 -60
rect 50 -400 130 -370
rect 50 -460 60 -400
rect 120 -460 130 -400
rect 50 -468 130 -460
rect 340 -400 420 -390
rect 340 -460 350 -400
rect 410 -460 420 -400
rect 340 -470 420 -460
rect 1370 -400 1450 -120
rect 1540 -60 1620 130
rect 2020 141 2100 200
rect 2080 80 2100 141
rect 2020 69 2100 80
rect 2850 100 2930 210
rect 3040 270 3140 280
rect 3040 190 3050 270
rect 3130 190 3140 270
rect 3410 270 3490 440
rect 3960 430 4040 450
rect 3960 370 3970 430
rect 4030 370 4040 430
rect 3780 340 3860 350
rect 3780 280 3790 340
rect 3850 280 3860 340
rect 3780 270 3860 280
rect 3960 270 4040 370
rect 4720 420 4800 430
rect 4720 360 4730 420
rect 4790 360 4800 420
rect 5490 400 5510 460
rect 4720 270 4800 360
rect 5070 350 5150 360
rect 5070 290 5080 350
rect 5140 290 5150 350
rect 5070 280 5150 290
rect 5490 280 5570 400
rect 6150 450 6300 480
rect 6150 390 6220 450
rect 6280 390 6300 450
rect 6150 370 6300 390
rect 5860 310 5940 320
rect 3040 180 3140 190
rect 3280 250 3360 260
rect 3280 190 3290 250
rect 3350 190 3360 250
rect 3410 210 3420 270
rect 3480 210 3490 270
rect 3410 200 3490 210
rect 3960 210 3970 270
rect 4030 210 4040 270
rect 3960 200 4040 210
rect 4160 250 4240 260
rect 2850 40 2860 100
rect 2920 40 2930 100
rect 2850 20 2930 40
rect 3280 100 3360 190
rect 3280 40 3290 100
rect 3350 40 3360 100
rect 3280 20 3360 40
rect 4160 190 4170 250
rect 4230 211 4240 250
rect 4360 250 4440 260
rect 4230 190 4241 211
rect 4160 121 4241 190
rect 4160 60 4170 121
rect 4230 60 4241 121
rect 4160 39 4241 60
rect 4360 190 4370 250
rect 4430 190 4440 250
rect 4700 210 4720 270
rect 4780 210 4800 270
rect 4700 200 4800 210
rect 4839 260 4920 269
rect 1540 -120 1550 -60
rect 1610 -120 1620 -60
rect 1540 -130 1620 -120
rect 4170 -30 4250 -20
rect 4170 -90 4180 -30
rect 4240 -90 4250 -30
rect 1490 -210 1570 -200
rect 1490 -270 1500 -210
rect 1560 -270 1570 -210
rect 3960 -220 4040 -210
rect 1490 -280 1570 -270
rect 2820 -230 2920 -220
rect 1500 -380 1560 -280
rect 2820 -310 2830 -230
rect 2910 -240 2920 -230
rect 2910 -310 2930 -240
rect 3960 -280 3970 -220
rect 3960 -290 4040 -280
rect 2820 -320 2930 -310
rect 1500 -390 1570 -380
rect 2850 -390 2930 -320
rect 1370 -460 1380 -400
rect 1440 -460 1450 -400
rect 1370 -470 1450 -460
rect 1490 -400 1570 -390
rect 1490 -460 1500 -400
rect 1560 -460 1570 -400
rect 1490 -470 1570 -460
rect 1630 -400 1710 -390
rect 1630 -460 1640 -400
rect 1700 -460 1710 -400
rect 2850 -450 2860 -390
rect 2920 -450 2930 -390
rect 2850 -460 2930 -450
rect 3120 -390 3220 -380
rect 1630 -470 1710 -460
rect 3120 -470 3130 -390
rect 3210 -470 3220 -390
rect 4170 -400 4250 -90
rect 4360 -30 4440 190
rect 4839 199 4850 260
rect 4910 199 4920 260
rect 5490 220 5500 280
rect 5560 220 5570 280
rect 5490 210 5570 220
rect 5670 270 5750 280
rect 5670 210 5680 270
rect 5740 210 5750 270
rect 5860 250 5870 310
rect 5930 250 5940 310
rect 6220 260 6300 370
rect 6780 450 6860 470
rect 6780 390 6790 450
rect 6850 390 6860 450
rect 6580 350 6660 360
rect 6580 290 6590 350
rect 6650 290 6660 350
rect 6580 280 6660 290
rect 6780 260 6860 390
rect 7520 440 7600 470
rect 7520 380 7530 440
rect 7590 380 7600 440
rect 7520 270 7600 380
rect 5860 240 5940 250
rect 6190 250 6330 260
rect 4839 140 4920 199
rect 4810 119 4920 140
rect 4810 60 4840 119
rect 4900 60 4920 119
rect 4810 40 4920 60
rect 5670 130 5750 210
rect 6190 190 6220 250
rect 6280 190 6330 250
rect 6190 170 6330 190
rect 6360 250 6440 260
rect 6360 190 6370 250
rect 6430 190 6440 250
rect 6780 200 6790 260
rect 6850 200 6860 260
rect 6780 190 6860 200
rect 6980 260 7059 270
rect 6980 200 6990 260
rect 7050 200 7059 260
rect 6360 130 6440 190
rect 5670 120 5790 130
rect 5670 60 5690 120
rect 5750 60 5790 120
rect 5280 40 5370 50
rect 4810 39 4840 40
rect 4360 -90 4370 -30
rect 4430 -90 4440 -30
rect 4360 -100 4440 -90
rect 5280 -30 5290 40
rect 5360 -30 5370 40
rect 5670 30 5790 60
rect 6339 100 6440 130
rect 6339 40 6370 100
rect 6430 40 6440 100
rect 6339 30 6440 40
rect 6980 90 7059 200
rect 7170 250 7250 260
rect 7170 190 7180 250
rect 7240 190 7250 250
rect 7170 180 7250 190
rect 7399 250 7480 260
rect 7399 190 7410 250
rect 7470 190 7480 250
rect 7520 210 7530 270
rect 7590 210 7600 270
rect 7900 330 7980 340
rect 7900 270 7910 330
rect 7970 270 7980 330
rect 7900 260 7980 270
rect 7520 200 7600 210
rect 7399 170 7480 190
rect 7400 120 7480 170
rect 6980 30 6990 90
rect 7050 30 7059 90
rect 6980 20 7059 30
rect 7380 100 7490 120
rect 7380 40 7410 100
rect 7470 40 7490 100
rect 7380 20 7490 40
rect 4170 -460 4180 -400
rect 4240 -460 4250 -400
rect 4170 -470 4250 -460
rect 4430 -400 4510 -390
rect 4430 -460 4440 -400
rect 4430 -470 4510 -460
rect 3120 -480 3220 -470
rect 2650 -510 2730 -498
rect 250 -520 340 -510
rect 250 -580 260 -520
rect 320 -570 340 -520
rect 250 -630 270 -580
rect 330 -630 340 -570
rect 1160 -520 1240 -510
rect 1160 -620 1170 -520
rect 1230 -620 1240 -520
rect 1160 -630 1240 -620
rect 2650 -570 2660 -510
rect 2720 -570 2730 -510
rect 250 -640 340 -630
rect 2650 -710 2730 -570
rect 3030 -520 3110 -510
rect 3030 -620 3040 -520
rect 3100 -620 3110 -520
rect 4320 -520 4400 -510
rect 4320 -580 4330 -520
rect 4390 -580 4400 -520
rect 2650 -770 2660 -710
rect 2720 -770 2730 -710
rect 2650 -780 2730 -770
rect 4320 -710 4400 -580
rect 4320 -770 4330 -710
rect 4390 -770 4400 -710
rect 820 -910 900 -870
rect 2020 -910 2120 -890
rect 430 -920 900 -910
rect -70 -950 10 -940
rect -70 -1010 -60 -950
rect 0 -1010 10 -950
rect 430 -980 440 -920
rect 500 -980 830 -920
rect 890 -980 900 -920
rect 430 -990 900 -980
rect 1720 -920 2040 -910
rect 1720 -980 1729 -920
rect 1789 -970 2040 -920
rect 2100 -970 2120 -910
rect 1789 -980 2120 -970
rect 1720 -990 2120 -980
rect 2720 -900 2820 -890
rect 2720 -980 2730 -900
rect 2810 -980 2820 -900
rect 2720 -990 2820 -980
rect -70 -1080 10 -1010
rect -70 -1140 -60 -1080
rect 0 -1140 10 -1080
rect -70 -1150 10 -1140
rect 50 -1080 130 -1070
rect 1339 -1080 1419 -1070
rect 50 -1180 60 -1080
rect 120 -1180 130 -1080
rect 50 -1190 130 -1180
rect 1230 -1088 1310 -1080
rect 1230 -1150 1240 -1088
rect 1300 -1150 1310 -1088
rect 1339 -1140 1350 -1080
rect 1410 -1140 1419 -1080
rect 1339 -1150 1419 -1140
rect 2720 -1080 2800 -990
rect 3220 -1000 3690 -990
rect 2720 -1140 2730 -1080
rect 2790 -1140 2800 -1080
rect 2720 -1150 2800 -1140
rect 2830 -1060 2930 -1050
rect 2830 -1140 2840 -1060
rect 2920 -1140 2930 -1060
rect 3220 -1060 3230 -1000
rect 3290 -1060 3690 -1000
rect 4320 -1060 4400 -770
rect 5280 -630 5370 -30
rect 5480 -80 5560 -70
rect 5480 -140 5490 -80
rect 5550 -140 5560 -80
rect 5480 -170 5560 -140
rect 7110 -80 7200 -70
rect 7110 -140 7120 -80
rect 7180 -140 7200 -80
rect 7110 -170 7200 -140
rect 5480 -330 5550 -170
rect 5800 -220 5880 -210
rect 5800 -280 5810 -220
rect 5870 -280 5880 -220
rect 5480 -340 5560 -330
rect 5480 -400 5490 -340
rect 5550 -400 5560 -340
rect 5480 -410 5560 -400
rect 5670 -390 5750 -380
rect 5280 -700 5290 -630
rect 5360 -700 5370 -630
rect 5670 -450 5680 -390
rect 5740 -450 5750 -390
rect 3220 -1070 3690 -1060
rect 3610 -1130 3620 -1070
rect 3680 -1130 3690 -1070
rect 3610 -1140 3690 -1130
rect 4020 -1070 4100 -1060
rect 4020 -1130 4030 -1070
rect 4090 -1130 4100 -1070
rect 2830 -1150 2930 -1140
rect 1230 -1160 1310 -1150
rect 1230 -1220 1290 -1160
rect 4020 -1210 4100 -1130
rect 4150 -1070 4400 -1060
rect 4520 -1000 4840 -990
rect 4520 -1060 4530 -1000
rect 4590 -1060 4770 -1000
rect 4830 -1060 4840 -1000
rect 4520 -1070 4840 -1060
rect 4150 -1130 4160 -1070
rect 4220 -1130 4400 -1070
rect 4150 -1140 4400 -1130
rect 4010 -1220 4110 -1210
rect 1230 -1240 1310 -1220
rect 1230 -1250 1330 -1240
rect 1230 -1330 1240 -1250
rect 1320 -1330 1330 -1250
rect 4010 -1300 4020 -1220
rect 4100 -1300 4110 -1220
rect 4010 -1310 4110 -1300
rect 5280 -1300 5370 -700
rect 5540 -660 5620 -650
rect 5540 -720 5550 -660
rect 5610 -720 5620 -660
rect 5540 -1080 5620 -720
rect 5670 -870 5750 -450
rect 5800 -400 5880 -280
rect 6990 -250 7070 -240
rect 6990 -310 7000 -250
rect 7060 -310 7070 -250
rect 5800 -460 5810 -400
rect 5870 -460 5880 -400
rect 5800 -660 5880 -460
rect 5940 -399 6020 -390
rect 5940 -460 5950 -399
rect 6010 -460 6020 -399
rect 5940 -470 6020 -460
rect 6990 -400 7070 -310
rect 6990 -460 7000 -400
rect 7060 -460 7070 -400
rect 6990 -470 7070 -460
rect 7120 -400 7200 -170
rect 8100 -100 8190 510
rect 8290 500 8380 510
rect 8290 440 8300 500
rect 8360 440 8380 500
rect 9030 500 9130 510
rect 8290 290 8380 440
rect 8290 230 8300 290
rect 8360 230 8380 290
rect 8650 450 8740 460
rect 8650 380 8660 450
rect 8730 380 8740 450
rect 9030 420 9040 500
rect 9120 420 9130 500
rect 9030 410 9130 420
rect 8650 370 8740 380
rect 8290 210 8380 230
rect 8500 260 8580 270
rect 8500 200 8510 260
rect 8570 200 8580 260
rect 8500 180 8580 200
rect 8480 130 8580 180
rect 8480 70 8500 130
rect 8560 70 8580 130
rect 8480 50 8580 70
rect 8100 -170 8110 -100
rect 8180 -170 8190 -100
rect 7120 -460 7130 -400
rect 7190 -460 7200 -400
rect 7120 -470 7200 -460
rect 7260 -400 7340 -390
rect 7260 -460 7270 -400
rect 7330 -460 7340 -400
rect 7260 -470 7340 -460
rect 6780 -520 6860 -510
rect 6780 -610 6790 -520
rect 6850 -610 6860 -520
rect 5800 -720 5810 -660
rect 5870 -720 5880 -660
rect 5800 -730 5880 -720
rect 8100 -770 8190 -170
rect 8310 -40 8390 -30
rect 8310 -100 8320 -40
rect 8380 -100 8390 -40
rect 8310 -230 8390 -100
rect 8310 -290 8320 -230
rect 8380 -290 8390 -230
rect 8310 -300 8390 -290
rect 8520 -190 8600 -180
rect 8520 -250 8530 -190
rect 8590 -250 8600 -190
rect 8520 -400 8600 -250
rect 8650 -190 8730 370
rect 9050 260 9130 410
rect 9440 340 9520 350
rect 9440 280 9450 340
rect 9510 280 9520 340
rect 9050 200 9060 260
rect 9120 200 9130 260
rect 9050 190 9130 200
rect 9210 260 9310 280
rect 9440 270 9520 280
rect 9210 200 9220 260
rect 9280 200 9310 260
rect 9210 190 9310 200
rect 9210 160 9290 190
rect 9190 130 9290 160
rect 9190 70 9210 130
rect 9270 70 9290 130
rect 9190 50 9290 70
rect 8650 -250 8660 -190
rect 8720 -250 8730 -190
rect 8650 -260 8730 -250
rect 8520 -460 8530 -400
rect 8590 -460 8600 -400
rect 8520 -470 8600 -460
rect 8780 -330 8860 -320
rect 8780 -390 8790 -330
rect 8850 -390 8860 -330
rect 8780 -410 8860 -390
rect 8780 -470 8790 -410
rect 8850 -470 8860 -410
rect 8780 -480 8860 -470
rect 8670 -510 8750 -500
rect 8100 -840 8110 -770
rect 8180 -840 8190 -770
rect 8100 -860 8190 -840
rect 8370 -550 8450 -540
rect 8370 -610 8380 -550
rect 8440 -610 8450 -550
rect 8670 -570 8680 -510
rect 8740 -570 8750 -510
rect 8670 -580 8750 -570
rect 5670 -930 5680 -870
rect 5740 -930 5750 -870
rect 6360 -900 6460 -880
rect 5670 -940 5750 -930
rect 6030 -910 6460 -900
rect 6030 -970 6050 -910
rect 6110 -970 6390 -910
rect 6450 -970 6460 -910
rect 6030 -980 6460 -970
rect 6850 -910 6930 -900
rect 6850 -970 6860 -910
rect 6920 -970 6930 -910
rect 5540 -1140 5550 -1080
rect 5610 -1140 5620 -1080
rect 5670 -1070 5750 -1060
rect 5670 -1130 5680 -1070
rect 5740 -1130 5750 -1070
rect 5670 -1140 5750 -1130
rect 6850 -1080 6930 -970
rect 8370 -1010 8450 -610
rect 8370 -1070 8380 -1010
rect 8440 -1070 8450 -1010
rect 8870 -1000 9120 -990
rect 8870 -1060 8880 -1000
rect 8940 -1060 9050 -1000
rect 9110 -1060 9120 -1000
rect 6850 -1140 6860 -1080
rect 6920 -1140 6930 -1080
rect 5540 -1150 5620 -1140
rect 6850 -1150 6930 -1140
rect 6970 -1080 7050 -1070
rect 8370 -1080 8450 -1070
rect 8490 -1070 8570 -1060
rect 8870 -1070 9120 -1060
rect 6970 -1140 6980 -1080
rect 7040 -1140 7050 -1080
rect 6970 -1150 7050 -1140
rect 8490 -1130 8500 -1070
rect 8560 -1130 8570 -1070
rect 7280 -1170 7800 -1160
rect 7280 -1230 7290 -1170
rect 7350 -1230 7730 -1170
rect 7790 -1230 7800 -1170
rect 7280 -1240 7800 -1230
rect 8490 -1210 8570 -1130
rect 8490 -1270 8500 -1210
rect 8560 -1270 8570 -1210
rect 8490 -1280 8570 -1270
rect 1230 -1340 1330 -1330
rect 5280 -1370 5290 -1300
rect 5360 -1370 5370 -1300
rect 5280 -1390 5370 -1370
<< via2 >>
rect -110 380 -50 440
rect 610 380 670 440
rect 70 100 130 160
rect 1160 380 1220 440
rect 990 270 1050 330
rect 1050 270 1060 330
rect 1910 370 1970 430
rect 2690 440 2750 500
rect 2280 280 2340 340
rect 3420 440 3480 500
rect 500 100 560 160
rect 1360 90 1420 150
rect 60 -50 120 10
rect 240 -50 300 10
rect -120 -280 -60 -220
rect 1380 -120 1440 -60
rect 350 -460 410 -400
rect 2020 80 2080 141
rect 3050 260 3130 270
rect 3050 200 3060 260
rect 3060 200 3120 260
rect 3120 200 3130 260
rect 3050 190 3130 200
rect 3970 370 4030 430
rect 3790 280 3850 340
rect 4730 360 4790 420
rect 5510 400 5570 460
rect 5080 290 5140 349
rect 6220 390 6280 450
rect 2860 40 2920 100
rect 3290 40 3350 100
rect 4170 60 4230 121
rect 1550 -120 1610 -60
rect 4180 -90 4240 -30
rect 1500 -270 1560 -210
rect 2830 -310 2910 -230
rect 3970 -280 4030 -220
rect 4030 -280 4040 -220
rect 1640 -460 1700 -400
rect 3130 -400 3210 -390
rect 3130 -460 3140 -400
rect 3140 -460 3200 -400
rect 3200 -460 3210 -400
rect 3130 -470 3210 -460
rect 5870 250 5930 310
rect 6790 390 6850 450
rect 6590 290 6650 350
rect 7530 380 7590 440
rect 4840 60 4900 119
rect 5690 60 5750 120
rect 4370 -90 4430 -30
rect 6370 40 6430 100
rect 7180 190 7240 250
rect 7910 270 7970 330
rect 6990 30 7050 90
rect 7410 40 7470 100
rect 4440 -460 4500 -400
rect 4500 -460 4510 -400
rect 270 -580 320 -570
rect 320 -580 330 -570
rect 270 -630 330 -580
rect 1170 -580 1230 -560
rect 1170 -620 1230 -580
rect 3040 -580 3100 -560
rect 3040 -620 3100 -580
rect 2660 -770 2720 -710
rect 4330 -770 4390 -710
rect -60 -1010 0 -950
rect 830 -980 890 -920
rect 2040 -970 2100 -910
rect 2730 -980 2810 -900
rect 60 -1141 120 -1120
rect 60 -1180 120 -1141
rect 1350 -1140 1410 -1080
rect 2840 -1070 2920 -1060
rect 2840 -1130 2850 -1070
rect 2850 -1130 2910 -1070
rect 2910 -1130 2920 -1070
rect 2840 -1140 2920 -1130
rect 5490 -140 5550 -80
rect 7120 -140 7180 -80
rect 5810 -280 5870 -220
rect 3620 -1130 3680 -1070
rect 4770 -1060 4830 -1000
rect 1240 -1330 1320 -1250
rect 4020 -1300 4100 -1220
rect 5550 -720 5610 -660
rect 7000 -310 7060 -250
rect 5950 -460 6010 -400
rect 8300 440 8360 500
rect 9040 420 9120 500
rect 8500 70 8560 130
rect 7270 -460 7330 -400
rect 6790 -580 6850 -550
rect 6790 -610 6850 -580
rect 5810 -720 5870 -660
rect 8320 -100 8380 -40
rect 8530 -250 8590 -190
rect 9450 280 9510 340
rect 9210 70 9270 130
rect 8660 -250 8720 -190
rect 8790 -390 8850 -330
rect 8380 -610 8440 -550
rect 8680 -570 8740 -510
rect 5680 -930 5740 -870
rect 6390 -970 6450 -910
rect 6860 -970 6920 -910
rect 5680 -1130 5740 -1070
rect 9050 -1060 9110 -1000
rect 6980 -1140 7040 -1080
rect 7730 -1230 7790 -1170
rect 8500 -1270 8560 -1210
<< metal3 >>
rect 2670 520 3540 530
rect -130 450 690 460
rect -130 370 -120 450
rect -38 440 690 450
rect -38 380 610 440
rect 670 380 690 440
rect -38 370 690 380
rect -130 360 690 370
rect 1140 450 2050 460
rect 1140 370 1150 450
rect 1230 430 2050 450
rect 2670 440 2680 520
rect 2760 500 3540 520
rect 2760 440 3420 500
rect 3480 440 3540 500
rect 8290 500 9170 510
rect 5490 470 6352 480
rect 2670 430 3540 440
rect 3950 440 4140 450
rect 1230 370 1910 430
rect 1970 370 2050 430
rect 1140 360 2050 370
rect 3950 360 3960 440
rect 4040 430 4140 440
rect 4040 420 4820 430
rect 4040 360 4730 420
rect 4790 360 4820 420
rect 5490 390 5500 470
rect 5580 450 6352 470
rect 5580 390 6220 450
rect 6280 390 6352 450
rect 5490 380 6352 390
rect 6780 460 7640 470
rect 6780 380 6790 460
rect 6870 440 7640 460
rect 6870 380 7530 440
rect 7590 380 7640 440
rect 8290 420 8300 500
rect 8380 420 9040 500
rect 9120 420 9170 500
rect 8290 410 8640 420
rect 8750 410 9170 420
rect 6780 370 7640 380
rect 2260 350 2360 360
rect 970 340 1070 350
rect 970 260 980 340
rect 1060 260 1070 340
rect 2260 270 2270 350
rect 2350 270 2360 350
rect 3770 350 3870 360
rect 3950 350 4820 360
rect 5060 360 5160 370
rect 2260 260 2360 270
rect 3040 270 3140 280
rect 970 250 1070 260
rect 3040 190 3050 270
rect 3130 190 3140 270
rect 3770 270 3780 350
rect 3860 270 3870 350
rect 5060 280 5070 360
rect 5150 280 5160 360
rect 6570 360 6670 370
rect 5060 270 5160 280
rect 5860 310 6030 320
rect 3770 260 3870 270
rect 5860 250 5870 310
rect 5930 250 5940 310
rect 5860 240 5940 250
rect 5930 230 5940 240
rect 6020 230 6030 310
rect 6570 270 6580 360
rect 6660 270 6670 360
rect 9430 350 9530 360
rect 7890 340 7990 350
rect 7890 260 7900 340
rect 7980 260 7990 340
rect 9430 270 9440 350
rect 9520 270 9530 350
rect 9430 260 9530 270
rect 5930 220 6030 230
rect 7170 250 7650 260
rect 7890 250 7990 260
rect 3040 180 3140 190
rect 7170 190 7180 250
rect 7240 190 7560 250
rect 7170 180 7560 190
rect 60 170 570 180
rect 7550 170 7560 180
rect 7640 170 7650 250
rect 60 90 70 170
rect 140 160 570 170
rect 140 100 500 160
rect 560 100 570 160
rect 140 90 570 100
rect 60 80 570 90
rect 1340 160 2140 170
rect 7550 160 7650 170
rect 1340 80 1350 160
rect 1430 141 2140 160
rect 1430 80 2020 141
rect 2080 80 2140 141
rect 8490 140 9320 150
rect 4150 130 4930 140
rect 8570 130 9320 140
rect 1340 70 2140 80
rect 2840 110 3360 120
rect 2840 30 2850 110
rect 2930 100 3360 110
rect 2930 40 3290 100
rect 3350 40 3360 100
rect 4150 50 4160 130
rect 4240 119 4930 130
rect 4240 60 4840 119
rect 4900 60 4930 119
rect 4240 50 4930 60
rect 4150 40 4930 50
rect 5670 120 6450 130
rect 5670 40 5680 120
rect 5760 100 6450 120
rect 5760 40 6370 100
rect 6430 40 6450 100
rect 2930 30 3360 40
rect 5670 30 6450 40
rect 6980 110 7490 120
rect 6980 30 6990 110
rect 7070 100 7490 110
rect 7070 40 7410 100
rect 7470 40 7490 100
rect 8570 70 9210 130
rect 9270 70 9320 130
rect 8570 60 9320 70
rect 8490 50 9320 60
rect 7070 30 7490 40
rect 2840 20 3360 30
rect 6980 20 7490 30
rect 50 10 310 20
rect 50 -50 60 10
rect 120 -50 240 10
rect 300 -50 310 10
rect 4170 -30 4440 -20
rect 9020 -30 9120 -10
rect 9240 -20 9340 -10
rect 9240 -30 9250 -20
rect 50 -60 310 -50
rect 1370 -60 1620 -50
rect 180 -80 280 -60
rect 1370 -120 1380 -60
rect 1440 -120 1550 -60
rect 1610 -120 1620 -60
rect 4170 -90 4180 -30
rect 4240 -90 4370 -30
rect 4430 -90 4440 -30
rect 8310 -40 9250 -30
rect 4170 -100 4440 -90
rect 5480 -80 7430 -70
rect 1370 -130 1620 -120
rect 5480 -140 5490 -80
rect 5550 -140 7120 -80
rect 7180 -140 7340 -80
rect 5480 -150 7340 -140
rect 7330 -160 7340 -150
rect 7420 -160 7430 -80
rect 8310 -100 8320 -40
rect 8380 -100 9250 -40
rect 9330 -100 9340 -20
rect 8310 -110 9340 -100
rect 7330 -170 7430 -160
rect 8520 -190 8780 -180
rect -130 -210 1830 -200
rect -130 -220 1500 -210
rect -130 -280 -120 -220
rect -60 -270 1500 -220
rect 1560 -270 1740 -210
rect -60 -280 1740 -270
rect -130 -290 -50 -280
rect 1730 -290 1740 -280
rect 1820 -290 1830 -210
rect 3960 -220 5880 -210
rect 1730 -300 1830 -290
rect 2820 -230 2920 -220
rect 2820 -310 2830 -230
rect 2910 -240 2920 -230
rect 3030 -230 3130 -220
rect 3030 -240 3040 -230
rect 2910 -310 3040 -240
rect 3120 -310 3130 -230
rect 3960 -280 3970 -220
rect 4040 -280 5810 -220
rect 5870 -280 5880 -220
rect 7540 -230 7640 -220
rect 7540 -240 7550 -230
rect 3960 -290 5880 -280
rect 6990 -250 7550 -240
rect 2820 -320 3130 -310
rect 6990 -310 7000 -250
rect 7060 -310 7550 -250
rect 7630 -310 7640 -230
rect 8520 -250 8530 -190
rect 8590 -250 8660 -190
rect 8720 -250 8780 -190
rect 8520 -260 8780 -250
rect 6990 -320 7640 -310
rect 9420 -310 9520 -300
rect 9420 -320 9430 -310
rect 8780 -330 9430 -320
rect 2240 -380 2340 -370
rect 3760 -380 3860 -370
rect 2240 -390 2250 -380
rect 320 -400 420 -390
rect 320 -480 330 -400
rect 410 -480 420 -400
rect 1630 -400 2250 -390
rect 1630 -460 1640 -400
rect 1700 -460 2250 -400
rect 2330 -460 2340 -380
rect 1630 -470 2340 -460
rect 3120 -390 3220 -380
rect 3760 -390 3770 -380
rect 3120 -470 3130 -390
rect 3210 -460 3770 -390
rect 3850 -460 3860 -380
rect 5050 -380 5150 -370
rect 5050 -390 5060 -380
rect 3210 -470 3860 -460
rect 4430 -400 5060 -390
rect 4430 -460 4440 -400
rect 4510 -460 5060 -400
rect 5140 -460 5150 -380
rect 6570 -380 6670 -370
rect 6570 -390 6580 -380
rect 4430 -470 5150 -460
rect 5940 -400 6580 -390
rect 5940 -460 5950 -400
rect 6010 -460 6580 -400
rect 6660 -460 6670 -380
rect 7880 -380 7980 -370
rect 7880 -389 7890 -380
rect 7460 -390 7890 -389
rect 5940 -470 6670 -460
rect 7260 -400 7890 -390
rect 7260 -460 7270 -400
rect 7330 -460 7890 -400
rect 7970 -460 7980 -380
rect 8780 -390 8790 -330
rect 8850 -390 9430 -330
rect 9510 -390 9520 -310
rect 8780 -400 9520 -390
rect 7260 -470 7980 -460
rect 3120 -480 3220 -470
rect 320 -490 420 -480
rect 8670 -510 8750 -500
rect 8670 -540 8680 -510
rect 970 -560 1070 -540
rect 3020 -550 3120 -540
rect 250 -570 980 -560
rect 250 -630 270 -570
rect 330 -630 980 -570
rect 250 -640 980 -630
rect 1060 -640 1070 -560
rect 1160 -560 3030 -550
rect 1160 -620 1170 -560
rect 1230 -620 3030 -560
rect 3110 -620 3120 -550
rect 6780 -550 8680 -540
rect 6780 -610 6790 -550
rect 6850 -610 8380 -550
rect 8440 -570 8680 -550
rect 8740 -570 8750 -510
rect 8440 -610 8750 -570
rect 6780 -620 8750 -610
rect 1160 -630 3120 -620
rect 970 -650 1070 -640
rect 5540 -660 5880 -650
rect 2650 -710 4400 -700
rect 2650 -770 2660 -710
rect 2720 -770 4330 -710
rect 4390 -770 4400 -710
rect 5540 -720 5550 -660
rect 5610 -720 5810 -660
rect 5870 -720 5880 -660
rect 5540 -730 5880 -720
rect 2650 -780 4400 -770
rect 5920 -850 6020 -840
rect 5920 -860 5930 -850
rect 810 -870 910 -860
rect 320 -930 420 -920
rect 320 -940 330 -930
rect -70 -950 330 -940
rect -70 -1010 -60 -950
rect 0 -1010 330 -950
rect 410 -1010 420 -930
rect 810 -950 820 -870
rect 900 -950 910 -870
rect 5670 -870 5930 -860
rect 3760 -890 3860 -880
rect 810 -960 830 -950
rect 820 -980 830 -960
rect 890 -960 910 -950
rect 2020 -900 2120 -890
rect 890 -980 900 -960
rect 820 -990 900 -980
rect 2020 -980 2030 -900
rect 2110 -980 2120 -900
rect 2020 -990 2120 -980
rect 2720 -900 3770 -890
rect 2720 -980 2730 -900
rect 2810 -960 3770 -900
rect 3850 -960 3860 -890
rect 5670 -930 5680 -870
rect 5740 -930 5930 -870
rect 6010 -930 6020 -850
rect 2810 -970 3860 -960
rect 2810 -980 2820 -970
rect 4760 -980 4840 -930
rect 5670 -940 6020 -930
rect 6360 -890 6460 -880
rect 6360 -970 6370 -890
rect 6450 -970 6460 -890
rect 7870 -890 7970 -880
rect 7870 -900 7880 -890
rect 6360 -980 6460 -970
rect 6850 -910 7880 -900
rect 6850 -970 6860 -910
rect 6920 -970 7880 -910
rect 7960 -970 7970 -890
rect 6850 -980 7970 -970
rect 9020 -980 9120 -970
rect 2720 -990 2820 -980
rect 4750 -990 4850 -980
rect -70 -1020 420 -1010
rect 3010 -1050 3110 -1040
rect 1730 -1060 1830 -1050
rect 1730 -1070 1740 -1060
rect 1340 -1080 1740 -1070
rect 970 -1100 1070 -1090
rect 970 -1110 980 -1100
rect 49 -1120 980 -1110
rect 49 -1180 60 -1120
rect 120 -1180 980 -1120
rect 1060 -1180 1070 -1100
rect 1340 -1140 1350 -1080
rect 1410 -1140 1740 -1080
rect 1820 -1140 1830 -1060
rect 1340 -1150 1830 -1140
rect 2830 -1060 2930 -1050
rect 3010 -1060 3020 -1050
rect 2830 -1140 2840 -1060
rect 2920 -1130 3020 -1060
rect 3100 -1130 3110 -1050
rect 2920 -1140 3110 -1130
rect 3600 -1060 3700 -1050
rect 3600 -1140 3610 -1060
rect 3690 -1140 3700 -1060
rect 4750 -1070 4760 -990
rect 4840 -1070 4850 -990
rect 6570 -1050 6670 -1040
rect 6570 -1060 6580 -1050
rect 4750 -1080 4850 -1070
rect 5670 -1070 6580 -1060
rect 5670 -1130 5680 -1070
rect 5740 -1130 6580 -1070
rect 6660 -1130 6670 -1050
rect 7330 -1060 7430 -1050
rect 7330 -1070 7340 -1060
rect 5670 -1140 6670 -1130
rect 6970 -1080 7340 -1070
rect 6970 -1140 6980 -1080
rect 7040 -1140 7340 -1080
rect 7420 -1140 7430 -1060
rect 9020 -1060 9030 -980
rect 9110 -1060 9120 -980
rect 9020 -1070 9120 -1060
rect 2830 -1150 2930 -1140
rect 3600 -1150 3700 -1140
rect 6970 -1150 7430 -1140
rect 7700 -1150 7800 -1140
rect 49 -1190 1070 -1180
rect 2210 -1210 2330 -1200
rect 1230 -1240 1310 -1220
rect 2210 -1240 2240 -1210
rect 1230 -1250 2240 -1240
rect 1230 -1330 1240 -1250
rect 1320 -1290 2240 -1250
rect 2320 -1290 2330 -1210
rect 3610 -1220 3690 -1150
rect 5050 -1210 5150 -1200
rect 4010 -1220 4110 -1210
rect 5050 -1220 5060 -1210
rect 1320 -1300 2330 -1290
rect 4010 -1300 4020 -1220
rect 4100 -1290 5060 -1220
rect 5140 -1290 5150 -1210
rect 7700 -1230 7710 -1150
rect 7790 -1230 7800 -1150
rect 9410 -1190 9510 -1180
rect 9410 -1200 9420 -1190
rect 7700 -1240 7800 -1230
rect 8490 -1210 9420 -1200
rect 8490 -1270 8500 -1210
rect 8560 -1270 9420 -1210
rect 9500 -1270 9510 -1190
rect 8490 -1280 9510 -1270
rect 4100 -1300 5150 -1290
rect 1320 -1330 1330 -1300
rect 4010 -1310 4110 -1300
rect 1230 -1340 1330 -1330
<< via3 >>
rect -120 440 -38 450
rect -120 380 -110 440
rect -110 380 -50 440
rect -50 380 -38 440
rect -120 370 -38 380
rect 1150 440 1230 450
rect 1150 380 1160 440
rect 1160 380 1220 440
rect 1220 380 1230 440
rect 2680 500 2760 520
rect 2680 440 2690 500
rect 2690 440 2750 500
rect 2750 440 2760 500
rect 1150 370 1230 380
rect 3960 430 4040 440
rect 3960 370 3970 430
rect 3970 370 4030 430
rect 4030 370 4040 430
rect 3960 360 4040 370
rect 5500 460 5580 470
rect 5500 400 5510 460
rect 5510 400 5570 460
rect 5570 400 5580 460
rect 5500 390 5580 400
rect 6790 450 6870 460
rect 6790 390 6850 450
rect 6850 390 6870 450
rect 6790 380 6870 390
rect 8300 440 8360 500
rect 8360 440 8380 500
rect 8300 420 8380 440
rect 980 330 1060 340
rect 980 270 990 330
rect 990 270 1060 330
rect 980 260 1060 270
rect 2270 340 2350 350
rect 2270 280 2280 340
rect 2280 280 2340 340
rect 2340 280 2350 340
rect 2270 270 2350 280
rect 3050 190 3130 270
rect 3780 340 3860 350
rect 3780 280 3790 340
rect 3790 280 3850 340
rect 3850 280 3860 340
rect 3780 270 3860 280
rect 5070 349 5150 360
rect 5070 290 5080 349
rect 5080 290 5140 349
rect 5140 290 5150 349
rect 5070 280 5150 290
rect 5940 230 6020 310
rect 6580 350 6660 360
rect 6580 290 6590 350
rect 6590 290 6650 350
rect 6650 290 6660 350
rect 6580 270 6660 290
rect 7900 330 7980 340
rect 7900 270 7910 330
rect 7910 270 7970 330
rect 7970 270 7980 330
rect 7900 260 7980 270
rect 9440 340 9520 350
rect 9440 280 9450 340
rect 9450 280 9510 340
rect 9510 280 9520 340
rect 9440 270 9520 280
rect 7560 170 7640 250
rect 70 160 140 170
rect 70 100 130 160
rect 130 100 140 160
rect 70 90 140 100
rect 1350 150 1430 160
rect 1350 90 1360 150
rect 1360 90 1420 150
rect 1420 90 1430 150
rect 1350 80 1430 90
rect 8490 130 8570 140
rect 2850 100 2930 110
rect 2850 40 2860 100
rect 2860 40 2920 100
rect 2920 40 2930 100
rect 4160 121 4240 130
rect 4160 60 4170 121
rect 4170 60 4230 121
rect 4230 60 4240 121
rect 4160 50 4240 60
rect 5680 60 5690 120
rect 5690 60 5750 120
rect 5750 60 5760 120
rect 5680 40 5760 60
rect 2850 30 2930 40
rect 6990 90 7070 110
rect 6990 30 7050 90
rect 7050 30 7070 90
rect 8490 70 8500 130
rect 8500 70 8560 130
rect 8560 70 8570 130
rect 8490 60 8570 70
rect 7340 -160 7420 -80
rect 9250 -100 9330 -20
rect 1740 -290 1820 -210
rect 3040 -310 3120 -230
rect 7550 -310 7630 -230
rect 330 -460 350 -400
rect 350 -460 410 -400
rect 330 -480 410 -460
rect 2250 -460 2330 -380
rect 3770 -460 3850 -380
rect 5060 -460 5140 -380
rect 6580 -460 6660 -380
rect 7890 -460 7970 -380
rect 9430 -390 9510 -310
rect 980 -640 1060 -560
rect 3030 -560 3110 -550
rect 3030 -620 3040 -560
rect 3040 -620 3100 -560
rect 3100 -620 3110 -560
rect 330 -1010 410 -930
rect 820 -920 900 -870
rect 820 -950 830 -920
rect 830 -950 890 -920
rect 890 -950 900 -920
rect 2030 -910 2110 -900
rect 2030 -970 2040 -910
rect 2040 -970 2100 -910
rect 2100 -970 2110 -910
rect 2030 -980 2110 -970
rect 3770 -960 3850 -890
rect 5930 -930 6010 -850
rect 6370 -910 6450 -890
rect 6370 -970 6390 -910
rect 6390 -970 6450 -910
rect 7880 -970 7960 -890
rect 980 -1180 1060 -1100
rect 1740 -1140 1820 -1060
rect 3020 -1130 3100 -1050
rect 3610 -1070 3690 -1060
rect 3610 -1130 3620 -1070
rect 3620 -1130 3680 -1070
rect 3680 -1130 3690 -1070
rect 3610 -1140 3690 -1130
rect 4760 -1000 4840 -990
rect 4760 -1060 4770 -1000
rect 4770 -1060 4830 -1000
rect 4830 -1060 4840 -1000
rect 4760 -1070 4840 -1060
rect 6580 -1130 6660 -1050
rect 7340 -1140 7420 -1060
rect 9030 -1000 9110 -980
rect 9030 -1060 9050 -1000
rect 9050 -1060 9110 -1000
rect 2240 -1290 2320 -1210
rect 5060 -1290 5140 -1210
rect 7710 -1170 7790 -1150
rect 7710 -1230 7730 -1170
rect 7730 -1230 7790 -1170
rect 9420 -1270 9500 -1190
<< metal4 >>
rect -120 460 -40 640
rect -130 450 -30 460
rect -130 370 -120 450
rect -38 370 -30 450
rect -130 360 -30 370
rect 70 180 150 630
rect 60 170 150 180
rect 60 90 70 170
rect 140 90 150 170
rect 60 80 150 90
rect 320 -390 400 630
rect 320 -400 420 -390
rect 320 -480 330 -400
rect 410 -480 420 -400
rect 320 -490 420 -480
rect 330 -920 410 -490
rect 820 -860 900 630
rect 1150 460 1230 650
rect 1140 450 1240 460
rect 1140 370 1150 450
rect 1230 370 1240 450
rect 1140 360 1240 370
rect 970 340 1070 350
rect 970 260 980 340
rect 1060 260 1070 340
rect 970 250 1070 260
rect 980 -540 1060 250
rect 1350 170 1430 670
rect 1340 160 1440 170
rect 1340 80 1350 160
rect 1430 80 1440 160
rect 1340 70 1440 80
rect 1730 -210 1830 -200
rect 1730 -290 1740 -210
rect 1820 -290 1830 -210
rect 1730 -300 1830 -290
rect 970 -560 1070 -540
rect 970 -640 980 -560
rect 1060 -640 1070 -560
rect 970 -650 1070 -640
rect 810 -870 910 -860
rect 320 -930 420 -920
rect 320 -1010 330 -930
rect 410 -1010 420 -930
rect 810 -950 820 -870
rect 900 -950 910 -870
rect 810 -960 910 -950
rect 320 -1020 420 -1010
rect 980 -1090 1060 -650
rect 1750 -1050 1830 -300
rect 2040 -890 2120 630
rect 2680 530 2760 640
rect 2670 520 2770 530
rect 2670 440 2680 520
rect 2760 440 2770 520
rect 2670 430 2770 440
rect 2260 350 2360 360
rect 2260 270 2270 350
rect 2350 270 2360 350
rect 2260 260 2360 270
rect 2280 -370 2340 260
rect 2850 120 2930 640
rect 3040 270 3140 280
rect 3040 190 3050 270
rect 3130 190 3140 270
rect 3040 180 3140 190
rect 2840 110 2960 120
rect 2840 30 2850 110
rect 2930 30 2960 110
rect 2840 20 2960 30
rect 3050 -220 3130 180
rect 3030 -230 3130 -220
rect 3030 -310 3040 -230
rect 3120 -310 3130 -230
rect 3030 -320 3130 -310
rect 2240 -380 2340 -370
rect 2240 -460 2250 -380
rect 2330 -460 2340 -380
rect 2240 -470 2340 -460
rect 2020 -900 2120 -890
rect 2020 -980 2030 -900
rect 2110 -980 2120 -900
rect 2020 -990 2120 -980
rect 1730 -1060 1830 -1050
rect 970 -1100 1070 -1090
rect 970 -1180 980 -1100
rect 1060 -1180 1070 -1100
rect 1730 -1140 1740 -1060
rect 1820 -1140 1830 -1060
rect 1730 -1150 1830 -1140
rect 970 -1190 1070 -1180
rect 2250 -1200 2330 -470
rect 3020 -550 3120 -540
rect 3020 -620 3030 -550
rect 3110 -620 3120 -550
rect 3020 -630 3120 -620
rect 3030 -1040 3110 -630
rect 3010 -1050 3110 -1040
rect 3610 -1050 3690 620
rect 3960 450 4040 640
rect 3950 440 4060 450
rect 3950 360 3960 440
rect 4040 360 4060 440
rect 3770 350 3870 360
rect 3950 350 4060 360
rect 3770 270 3780 350
rect 3860 270 3870 350
rect 3770 260 3870 270
rect 3780 -370 3860 260
rect 4160 140 4240 640
rect 4150 130 4250 140
rect 4150 50 4160 130
rect 4240 50 4250 130
rect 4150 40 4250 50
rect 3760 -380 3860 -370
rect 3760 -460 3770 -380
rect 3850 -460 3860 -380
rect 3760 -470 3860 -460
rect 3780 -880 3860 -470
rect 3760 -890 3860 -880
rect 3760 -960 3770 -890
rect 3850 -960 3860 -890
rect 3760 -970 3860 -960
rect 4760 -980 4840 620
rect 5500 480 5580 640
rect 5490 470 5610 480
rect 5490 390 5500 470
rect 5580 390 5610 470
rect 5490 380 5610 390
rect 5060 360 5160 370
rect 5060 280 5070 360
rect 5150 280 5160 360
rect 5060 270 5160 280
rect 5070 -370 5150 270
rect 5680 130 5760 640
rect 5930 310 6030 320
rect 5930 230 5940 310
rect 6020 230 6030 310
rect 5930 220 6030 230
rect 5670 120 5780 130
rect 5670 40 5680 120
rect 5760 40 5780 120
rect 5670 30 5780 40
rect 5050 -380 5150 -370
rect 5050 -460 5060 -380
rect 5140 -460 5150 -380
rect 5050 -470 5150 -460
rect 4750 -990 4850 -980
rect 3010 -1130 3020 -1050
rect 3100 -1130 3110 -1050
rect 3010 -1140 3110 -1130
rect 3600 -1060 3700 -1050
rect 3600 -1140 3610 -1060
rect 3690 -1140 3700 -1060
rect 4750 -1070 4760 -990
rect 4840 -1070 4850 -990
rect 4750 -1080 4850 -1070
rect 3600 -1150 3700 -1140
rect 5070 -1200 5150 -470
rect 5940 -840 6020 220
rect 5920 -850 6020 -840
rect 5920 -930 5930 -850
rect 6010 -930 6020 -850
rect 6380 -880 6460 620
rect 6790 470 6870 670
rect 6780 460 6890 470
rect 6780 380 6790 460
rect 6870 380 6890 460
rect 6780 370 6890 380
rect 6570 360 6670 370
rect 6570 270 6580 360
rect 6660 270 6670 360
rect 6570 260 6670 270
rect 6590 -370 6670 260
rect 6990 120 7070 670
rect 7550 250 7650 260
rect 7550 170 7560 250
rect 7640 170 7650 250
rect 7550 160 7650 170
rect 6980 110 7089 120
rect 6980 30 6990 110
rect 7070 30 7089 110
rect 6980 20 7089 30
rect 7330 -80 7430 -70
rect 7330 -160 7340 -80
rect 7420 -160 7430 -80
rect 7330 -170 7430 -160
rect 6570 -380 6670 -370
rect 6570 -460 6580 -380
rect 6660 -460 6670 -380
rect 6570 -470 6670 -460
rect 5920 -940 6020 -930
rect 6360 -890 6460 -880
rect 6360 -970 6370 -890
rect 6450 -970 6460 -890
rect 6360 -980 6460 -970
rect 6590 -1040 6670 -470
rect 6570 -1050 6670 -1040
rect 7350 -1050 7430 -170
rect 7560 -220 7640 160
rect 7540 -230 7640 -220
rect 7540 -310 7550 -230
rect 7630 -310 7640 -230
rect 7540 -320 7640 -310
rect 6570 -1130 6580 -1050
rect 6660 -1130 6670 -1050
rect 6570 -1140 6670 -1130
rect 7330 -1060 7430 -1050
rect 7330 -1140 7340 -1060
rect 7420 -1140 7430 -1060
rect 7720 -1140 7800 640
rect 8300 510 8380 650
rect 8290 500 8430 510
rect 8290 420 8300 500
rect 8380 420 8430 500
rect 8290 410 8430 420
rect 7890 340 7990 350
rect 7890 260 7900 340
rect 7980 260 7990 340
rect 7890 250 7990 260
rect 7900 -370 7980 250
rect 8490 180 8570 650
rect 8480 140 8580 180
rect 8480 60 8490 140
rect 8570 60 8580 140
rect 8480 50 8580 60
rect 9040 -10 9120 620
rect 9260 -10 9340 620
rect 9430 350 9530 360
rect 9430 270 9440 350
rect 9520 270 9530 350
rect 9430 260 9530 270
rect 9020 -110 9120 -10
rect 9240 -20 9340 -10
rect 9240 -100 9250 -20
rect 9330 -100 9340 -20
rect 9240 -110 9340 -100
rect 7880 -380 7980 -370
rect 7880 -460 7890 -380
rect 7970 -460 7980 -380
rect 7880 -470 7980 -460
rect 7890 -880 7970 -470
rect 7870 -890 7970 -880
rect 7870 -970 7880 -890
rect 7960 -970 7970 -890
rect 9040 -970 9120 -110
rect 9440 -300 9520 260
rect 9420 -310 9520 -300
rect 9420 -390 9430 -310
rect 9510 -390 9520 -310
rect 9420 -400 9520 -390
rect 7870 -980 7970 -970
rect 9020 -980 9120 -970
rect 9020 -1060 9030 -980
rect 9110 -1060 9120 -980
rect 9020 -1070 9120 -1060
rect 7330 -1150 7430 -1140
rect 7700 -1150 7800 -1140
rect 2210 -1210 2330 -1200
rect 2210 -1290 2240 -1210
rect 2320 -1290 2330 -1210
rect 2210 -1300 2330 -1290
rect 5050 -1210 5150 -1200
rect 5050 -1290 5060 -1210
rect 5140 -1290 5150 -1210
rect 7700 -1230 7710 -1150
rect 7790 -1230 7800 -1150
rect 9430 -1180 9510 -400
rect 7700 -1240 7800 -1230
rect 9410 -1190 9510 -1180
rect 9410 -1270 9420 -1190
rect 9500 -1270 9510 -1190
rect 9410 -1280 9510 -1270
rect 5050 -1300 5150 -1290
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_0
timestamp 1747071801
transform 1 0 -132 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_1
timestamp 1747071801
transform 1 0 1162 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_2
timestamp 1747071801
transform 1 0 2658 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_3
timestamp 1747071801
transform 1 0 3954 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_4
timestamp 1747071801
transform 1 0 5478 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_5
timestamp 1747071801
transform 1 0 6788 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_6
timestamp 1747071801
transform 1 0 8310 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0
timestamp 1747071801
transform 1 0 -132 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_1
timestamp 1747071801
transform 1 0 1160 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_2
timestamp 1747071801
transform 1 0 2658 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_3
timestamp 1747071801
transform 1 0 3968 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_4
timestamp 1747071801
transform 1 0 5478 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_5
timestamp 1747071801
transform 1 0 6788 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_6
timestamp 1747071801
transform 1 0 8310 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0
timestamp 1747071801
transform 1 0 664 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1747071801
transform 1 0 1922 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_2
timestamp 1747071801
transform 1 0 9166 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_3
timestamp 1747071801
transform 1 0 3437 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_4
timestamp 1747071801
transform 1 0 4757 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_5
timestamp 1747071801
transform 1 0 6273 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_6
timestamp 1747071801
transform 1 0 7578 0 1 -1342
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_0
timestamp 1747071801
transform 1 0 518 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_1
timestamp 1747071801
transform 1 0 1804 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_2
timestamp 1747071801
transform 1 0 3306 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_3
timestamp 1747071801
transform 1 0 4600 0 1 -670
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_4
timestamp 1747071801
transform 1 0 6118 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_5
timestamp 1747071801
transform 1 0 7428 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_6
timestamp 1747071801
transform 1 0 8982 0 1 -668
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1747071801
transform 1 0 2448 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1747071801
transform 1 0 5278 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1747071801
transform 1 0 8100 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1747071801
transform 1 0 2448 0 1 -670
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1747071801
transform 1 0 2448 0 1 -1342
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1747071801
transform 1 0 5278 0 1 -668
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1747071801
transform 1 0 5278 0 1 -1342
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1747071801
transform 1 0 8100 0 1 -668
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1747071801
transform 1 0 8100 0 1 -1342
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0
timestamp 1747333433
transform 1 0 422 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1747333433
transform 1 0 1710 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_2
timestamp 1747333433
transform 1 0 3228 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_3
timestamp 1747333433
transform 1 0 4528 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_4
timestamp 1747333433
transform 1 0 6038 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_5
timestamp 1747333433
transform 1 0 7348 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_6
timestamp 1747333433
transform 1 0 8890 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_7
timestamp 1747333433
transform 1 0 -132 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_8
timestamp 1747333433
transform 1 0 1162 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_9
timestamp 1747333433
transform 1 0 2658 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_10
timestamp 1747333433
transform 1 0 3954 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_11
timestamp 1747333433
transform 1 0 5478 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_12
timestamp 1747333433
transform 1 0 6788 0 1 -1342
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_13
timestamp 1747333433
transform 1 0 8308 0 1 -1342
box -38 -48 682 592
<< labels >>
rlabel metal4 850 610 850 610 7 S1
port 4 w
rlabel metal4 2080 610 2080 610 7 S2
port 7 w
rlabel metal4 2720 610 2720 610 7 A3
port 8 w
rlabel metal4 2890 620 2890 620 7 B3
port 9 w
rlabel metal4 3650 610 3650 610 7 S3
port 10 w
rlabel metal4 4000 620 4000 620 7 A4
port 11 w
rlabel metal4 4200 620 4200 620 7 B4
port 12 w
rlabel metal4 4800 600 4800 600 7 S4
port 13 w
rlabel metal4 5540 620 5540 620 7 A5
port 14 w
rlabel metal4 5710 620 5710 620 7 B5
port 15 w
rlabel metal4 6410 600 6410 600 7 S5
port 16 w
rlabel metal4 6820 640 6820 640 7 A6
port 17 w
rlabel metal4 7020 630 7020 630 7 B6
port 18 w
rlabel metal4 7750 610 7750 610 7 S6
port 19 w
rlabel metal4 8330 620 8330 620 7 A7
port 20 w
rlabel metal4 8530 620 8530 620 7 B7
port 21 w
rlabel metal4 9080 610 9080 610 7 S7
port 22 w
rlabel metal4 9290 610 9290 610 7 CO
port 23 w
rlabel metal1 s 40 540 40 540 7 VDD_1
port 24 w
rlabel metal1 s 40 -1340 40 -1340 7 GND_3
port 29 w
rlabel metal4 -90 620 -90 620 7 A1
port 1 w
rlabel metal4 110 610 110 610 7 B1
port 2 w
rlabel metal4 370 610 370 610 7 CI
port 3 w
rlabel metal4 1180 620 1180 620 7 A2
port 5 w
rlabel metal4 1390 620 1390 620 7 B2
port 6 w
<< end >>
