magic
tech sky130A
timestamp 1747161529
<< metal1 >>
rect 3085 20120 3115 20150
rect 3085 20055 3115 20085
rect 3085 19785 3115 19815
rect 3085 19715 3115 19745
<< via1 >>
rect 3020 20390 3050 20420
rect 3085 19450 3115 19480
<< metal2 >>
rect 2945 20420 3055 20430
rect 2945 20390 2950 20420
rect 2980 20390 3020 20420
rect 3050 20390 3055 20420
rect 2945 20380 3055 20390
rect 3080 19480 3120 19490
rect 3080 19450 3085 19480
rect 3115 19450 3120 19480
rect 3080 19440 3120 19450
<< via2 >>
rect 2950 20390 2980 20420
rect 3085 19450 3115 19480
<< metal3 >>
rect 2710 22430 14720 22435
rect 2710 22390 2715 22430
rect 2755 22390 3065 22430
rect 3105 22390 3240 22430
rect 3280 22390 3340 22430
rect 3380 22390 3615 22430
rect 3655 22390 3890 22430
rect 3930 22390 4165 22430
rect 4205 22390 4440 22430
rect 4480 22390 4715 22430
rect 4755 22390 4990 22430
rect 5030 22390 5270 22430
rect 5310 22390 5545 22430
rect 5585 22390 5820 22430
rect 5860 22390 6100 22430
rect 6140 22390 6375 22430
rect 6415 22390 6650 22430
rect 6690 22390 6925 22430
rect 6965 22390 7205 22430
rect 7245 22390 14720 22430
rect 2710 22385 14720 22390
rect 3060 22340 14720 22345
rect 3060 22300 4885 22340
rect 4925 22300 8860 22340
rect 8900 22300 14720 22340
rect 3060 22295 14720 22300
rect 3060 22250 14720 22255
rect 3060 22210 4505 22250
rect 4545 22210 12445 22250
rect 12485 22210 14720 22250
rect 3060 22205 14720 22210
rect 3060 22160 14720 22165
rect 3060 22120 4420 22160
rect 4460 22120 12725 22160
rect 12765 22120 14720 22160
rect 3060 22115 14720 22120
rect 3060 22070 14720 22075
rect 3060 22030 4100 22070
rect 4140 22030 9135 22070
rect 9175 22030 14720 22070
rect 3060 22025 14720 22030
rect 400 21980 2760 21985
rect 400 21940 405 21980
rect 445 21940 470 21980
rect 510 21940 535 21980
rect 575 21940 2715 21980
rect 2755 21940 2760 21980
rect 400 21935 2760 21940
rect 3060 21980 14720 21985
rect 3060 21940 3755 21980
rect 3795 21940 13000 21980
rect 13040 21940 14720 21980
rect 3060 21935 14720 21940
rect 3060 21890 14720 21895
rect 3060 21850 3655 21890
rect 3695 21850 13275 21890
rect 13315 21850 14720 21890
rect 3060 21845 14720 21850
rect 3060 21800 14720 21805
rect 3060 21760 7480 21800
rect 7520 21760 7710 21800
rect 7750 21760 14720 21800
rect 3060 21755 14720 21760
rect 3060 21710 14720 21715
rect 3060 21670 7600 21710
rect 7640 21670 7875 21710
rect 7915 21670 14720 21710
rect 3060 21665 14385 21670
rect 3015 21620 14720 21625
rect 3015 21580 7325 21620
rect 7365 21580 10240 21620
rect 10280 21580 14720 21620
rect 3015 21575 14720 21580
rect 3015 21530 14720 21535
rect 3015 21490 7230 21530
rect 7270 21490 10515 21530
rect 10555 21490 14720 21530
rect 3015 21485 14720 21490
rect 3015 21440 14720 21445
rect 3015 21400 6940 21440
rect 6980 21400 8025 21440
rect 8065 21400 14720 21440
rect 3015 21395 14720 21400
rect 3015 21350 14720 21355
rect 3015 21310 6575 21350
rect 6615 21310 10790 21350
rect 10830 21310 14720 21350
rect 3015 21305 14720 21310
rect 3015 21260 14720 21265
rect 3015 21220 6475 21260
rect 6515 21220 11065 21260
rect 11105 21220 14720 21260
rect 3015 21215 14720 21220
rect 6265 21175 6315 21180
rect 8300 21175 8350 21180
rect 3015 21135 6270 21175
rect 6310 21135 8305 21175
rect 8345 21135 14720 21175
rect 6265 21130 6315 21135
rect 8300 21130 8350 21135
rect 5915 21095 5965 21100
rect 11340 21095 11390 21100
rect 3015 21055 5920 21095
rect 5960 21055 11345 21095
rect 11385 21055 14720 21095
rect 5915 21050 5965 21055
rect 11340 21050 11390 21055
rect 5825 21015 5875 21020
rect 11615 21015 11665 21020
rect 3015 20975 5830 21015
rect 5870 20975 11620 21015
rect 11660 20975 14720 21015
rect 5825 20970 5875 20975
rect 11615 20970 11665 20975
rect 5455 20935 5505 20940
rect 8580 20935 8630 20940
rect 3015 20895 5460 20935
rect 5500 20895 8585 20935
rect 8625 20895 14720 20935
rect 5455 20890 5505 20895
rect 8580 20890 8630 20895
rect 5155 20855 5205 20860
rect 11890 20855 11940 20860
rect 3015 20815 5160 20855
rect 5200 20815 11895 20855
rect 11935 20815 14720 20855
rect 5155 20810 5205 20815
rect 11890 20810 11940 20815
rect 5055 20775 5105 20780
rect 12165 20775 12215 20780
rect 3015 20735 5060 20775
rect 5100 20735 12170 20775
rect 12210 20735 14720 20775
rect 5055 20730 5105 20735
rect 12165 20730 12215 20735
rect 3485 20695 3535 20700
rect 3015 20655 3490 20695
rect 3530 20655 9410 20695
rect 9450 20655 14720 20695
rect 3485 20650 3535 20655
rect 3110 20615 3160 20620
rect 13540 20615 13590 20620
rect 3015 20575 3115 20615
rect 3155 20575 13545 20615
rect 13585 20575 14720 20615
rect 3110 20570 3160 20575
rect 13540 20570 13590 20575
rect 3015 20535 3065 20540
rect 13820 20535 13870 20540
rect 3015 20495 3020 20535
rect 3060 20495 13825 20535
rect 13865 20495 14720 20535
rect 3015 20490 3065 20495
rect 13820 20490 13870 20495
rect 100 20425 2985 20430
rect 100 20385 110 20425
rect 150 20385 175 20425
rect 215 20385 240 20425
rect 280 20420 2985 20425
rect 280 20390 2950 20420
rect 2980 20390 2985 20420
rect 280 20385 2985 20390
rect 100 20380 2985 20385
rect 400 19485 3120 19490
rect 400 19445 410 19485
rect 450 19445 475 19485
rect 515 19445 540 19485
rect 580 19480 3120 19485
rect 580 19450 3085 19480
rect 3115 19450 3120 19480
rect 580 19445 3120 19450
rect 400 19440 3120 19445
<< via3 >>
rect 2715 22390 2755 22430
rect 3065 22390 3105 22430
rect 3240 22390 3280 22430
rect 3340 22390 3380 22430
rect 3615 22390 3655 22430
rect 3890 22390 3930 22430
rect 4165 22390 4205 22430
rect 4440 22390 4480 22430
rect 4715 22390 4755 22430
rect 4990 22390 5030 22430
rect 5270 22390 5310 22430
rect 5545 22390 5585 22430
rect 5820 22390 5860 22430
rect 6100 22390 6140 22430
rect 6375 22390 6415 22430
rect 6650 22390 6690 22430
rect 6925 22390 6965 22430
rect 7205 22390 7245 22430
rect 4885 22300 4925 22340
rect 8860 22300 8900 22340
rect 4505 22210 4545 22250
rect 12445 22210 12485 22250
rect 4420 22120 4460 22160
rect 12725 22120 12765 22160
rect 4100 22030 4140 22070
rect 9135 22030 9175 22070
rect 405 21940 445 21980
rect 470 21940 510 21980
rect 535 21940 575 21980
rect 2715 21940 2755 21980
rect 3755 21940 3795 21980
rect 13000 21940 13040 21980
rect 3655 21850 3695 21890
rect 13275 21850 13315 21890
rect 7480 21760 7520 21800
rect 7710 21760 7750 21800
rect 7600 21670 7640 21710
rect 7875 21670 7915 21710
rect 7325 21580 7365 21620
rect 10240 21580 10280 21620
rect 7230 21490 7270 21530
rect 10515 21490 10555 21530
rect 6940 21400 6980 21440
rect 8025 21400 8065 21440
rect 6575 21310 6615 21350
rect 10790 21310 10830 21350
rect 6475 21220 6515 21260
rect 11065 21220 11105 21260
rect 6270 21135 6310 21175
rect 8305 21135 8345 21175
rect 5920 21055 5960 21095
rect 11345 21055 11385 21095
rect 5830 20975 5870 21015
rect 11620 20975 11660 21015
rect 5460 20895 5500 20935
rect 8585 20895 8625 20935
rect 5160 20815 5200 20855
rect 11895 20815 11935 20855
rect 5060 20735 5100 20775
rect 12170 20735 12210 20775
rect 3490 20655 3530 20695
rect 9410 20655 9450 20695
rect 3115 20575 3155 20615
rect 13545 20575 13585 20615
rect 3020 20495 3060 20535
rect 13825 20495 13865 20535
rect 110 20385 150 20425
rect 175 20385 215 20425
rect 240 20385 280 20425
rect 410 19445 450 19485
rect 475 19445 515 19485
rect 540 19445 580 19485
<< metal4 >>
rect 3067 22485 3097 22576
rect 3343 22485 3373 22576
rect 3619 22485 3649 22576
rect 3895 22485 3925 22576
rect 4171 22485 4201 22576
rect 4447 22485 4477 22576
rect 4723 22485 4753 22576
rect 4999 22485 5029 22576
rect 5275 22495 5305 22576
rect 3065 22435 3105 22485
rect 3340 22435 3380 22485
rect 3615 22435 3655 22485
rect 3890 22435 3930 22485
rect 4165 22435 4205 22485
rect 4440 22435 4480 22485
rect 4715 22435 4755 22485
rect 4990 22435 5030 22485
rect 5270 22435 5310 22495
rect 5551 22490 5581 22576
rect 5827 22490 5857 22576
rect 6103 22490 6133 22576
rect 6379 22495 6409 22576
rect 5545 22435 5585 22490
rect 5820 22435 5860 22490
rect 6100 22435 6140 22490
rect 6375 22435 6415 22495
rect 6655 22490 6685 22576
rect 6931 22505 6961 22576
rect 6650 22435 6690 22490
rect 6925 22435 6965 22505
rect 7207 22490 7237 22576
rect 7483 22490 7513 22576
rect 7759 22490 7789 22576
rect 8035 22550 8065 22576
rect 7205 22435 7245 22490
rect 2710 22430 2760 22435
rect 2710 22390 2715 22430
rect 2755 22390 2760 22430
rect 2710 22385 2760 22390
rect 3060 22430 3110 22435
rect 3060 22390 3065 22430
rect 3105 22390 3110 22430
rect 3060 22385 3110 22390
rect 3235 22430 3285 22435
rect 3235 22390 3240 22430
rect 3280 22390 3285 22430
rect 3235 22385 3285 22390
rect 3335 22430 3385 22435
rect 3335 22390 3340 22430
rect 3380 22390 3385 22430
rect 3335 22385 3385 22390
rect 3610 22430 3660 22435
rect 3610 22390 3615 22430
rect 3655 22390 3660 22430
rect 3610 22385 3660 22390
rect 3885 22430 3935 22435
rect 3885 22390 3890 22430
rect 3930 22390 3935 22430
rect 3885 22385 3935 22390
rect 4160 22430 4210 22435
rect 4160 22390 4165 22430
rect 4205 22390 4210 22430
rect 4160 22385 4210 22390
rect 4435 22430 4485 22435
rect 4435 22390 4440 22430
rect 4480 22390 4485 22430
rect 4435 22385 4485 22390
rect 4710 22430 4760 22435
rect 4710 22390 4715 22430
rect 4755 22390 4760 22430
rect 4710 22385 4760 22390
rect 4985 22430 5035 22435
rect 4985 22390 4990 22430
rect 5030 22390 5035 22430
rect 4985 22385 5035 22390
rect 5265 22430 5315 22435
rect 5265 22390 5270 22430
rect 5310 22390 5315 22430
rect 5265 22385 5315 22390
rect 5540 22430 5590 22435
rect 5540 22390 5545 22430
rect 5585 22390 5590 22430
rect 5540 22385 5590 22390
rect 5815 22430 5865 22435
rect 5815 22390 5820 22430
rect 5860 22390 5865 22430
rect 5815 22385 5865 22390
rect 6095 22430 6145 22435
rect 6095 22390 6100 22430
rect 6140 22390 6145 22430
rect 6095 22385 6145 22390
rect 6370 22430 6420 22435
rect 6370 22390 6375 22430
rect 6415 22390 6420 22430
rect 6370 22385 6420 22390
rect 6645 22430 6695 22435
rect 6645 22390 6650 22430
rect 6690 22390 6695 22430
rect 6645 22385 6695 22390
rect 6920 22430 6970 22435
rect 6920 22390 6925 22430
rect 6965 22390 6970 22430
rect 6920 22385 6970 22390
rect 7200 22430 7250 22435
rect 7200 22390 7205 22430
rect 7245 22390 7250 22430
rect 7200 22385 7250 22390
rect 100 20425 300 22076
rect 100 20385 110 20425
rect 150 20385 175 20425
rect 215 20385 240 20425
rect 280 20385 300 20425
rect 100 500 300 20385
rect 400 21980 600 22076
rect 2715 21985 2755 22385
rect 400 21940 405 21980
rect 445 21940 470 21980
rect 510 21940 535 21980
rect 575 21940 600 21980
rect 400 19485 600 21940
rect 2710 21980 2760 21985
rect 2710 21940 2715 21980
rect 2755 21940 2760 21980
rect 2710 21935 2760 21940
rect 3110 20615 3160 20620
rect 3110 20575 3115 20615
rect 3155 20575 3160 20615
rect 3110 20570 3160 20575
rect 3015 20535 3065 20540
rect 3015 20495 3020 20535
rect 3060 20495 3065 20535
rect 3015 20490 3065 20495
rect 3020 20445 3060 20490
rect 3115 20440 3155 20570
rect 3240 20445 3280 22385
rect 4880 22340 4930 22345
rect 4880 22300 4885 22340
rect 4925 22300 4930 22340
rect 4880 22295 4930 22300
rect 4500 22250 4550 22255
rect 4500 22210 4505 22250
rect 4545 22210 4550 22250
rect 4500 22205 4550 22210
rect 4415 22160 4465 22165
rect 4415 22120 4420 22160
rect 4460 22120 4465 22160
rect 4415 22115 4465 22120
rect 4095 22070 4145 22075
rect 4095 22030 4100 22070
rect 4140 22030 4145 22070
rect 4095 22025 4145 22030
rect 3750 21980 3800 21985
rect 3750 21940 3755 21980
rect 3795 21940 3800 21980
rect 3750 21935 3800 21940
rect 3650 21890 3700 21895
rect 3650 21850 3655 21890
rect 3695 21850 3700 21890
rect 3650 21845 3700 21850
rect 3485 20695 3535 20700
rect 3485 20655 3490 20695
rect 3530 20655 3535 20695
rect 3485 20650 3535 20655
rect 3490 20440 3530 20650
rect 3655 20445 3695 21845
rect 3755 20445 3795 21935
rect 4100 20440 4140 22025
rect 4420 20445 4460 22115
rect 4505 20445 4545 22205
rect 4885 20435 4925 22295
rect 7480 21805 7520 22490
rect 7755 22435 7795 22490
rect 7755 22385 7915 22435
rect 7475 21800 7525 21805
rect 7475 21760 7480 21800
rect 7520 21760 7525 21800
rect 7475 21755 7525 21760
rect 7705 21800 7755 21805
rect 7705 21760 7710 21800
rect 7750 21760 7755 21800
rect 7705 21755 7755 21760
rect 7595 21710 7645 21715
rect 7595 21670 7600 21710
rect 7640 21670 7645 21710
rect 7595 21665 7645 21670
rect 7320 21620 7370 21625
rect 7320 21580 7325 21620
rect 7365 21580 7370 21620
rect 7320 21575 7370 21580
rect 7225 21530 7275 21535
rect 7225 21490 7230 21530
rect 7270 21490 7275 21530
rect 7225 21485 7275 21490
rect 6935 21440 6985 21445
rect 6935 21400 6940 21440
rect 6980 21400 6985 21440
rect 6935 21395 6985 21400
rect 6570 21350 6620 21355
rect 6570 21310 6575 21350
rect 6615 21310 6620 21350
rect 6570 21305 6620 21310
rect 6470 21260 6520 21265
rect 6470 21220 6475 21260
rect 6515 21220 6520 21260
rect 6470 21215 6520 21220
rect 6265 21175 6315 21180
rect 6265 21135 6270 21175
rect 6310 21135 6315 21175
rect 6265 21130 6315 21135
rect 5915 21095 5965 21100
rect 5915 21055 5920 21095
rect 5960 21055 5965 21095
rect 5915 21050 5965 21055
rect 5825 21015 5875 21020
rect 5825 20975 5830 21015
rect 5870 20975 5875 21015
rect 5825 20970 5875 20975
rect 5455 20935 5505 20940
rect 5455 20895 5460 20935
rect 5500 20895 5505 20935
rect 5455 20890 5505 20895
rect 5155 20855 5205 20860
rect 5155 20815 5160 20855
rect 5200 20815 5205 20855
rect 5155 20810 5205 20815
rect 5055 20775 5105 20780
rect 5055 20735 5060 20775
rect 5100 20735 5105 20775
rect 5055 20730 5105 20735
rect 5060 20440 5100 20730
rect 5160 20445 5200 20810
rect 5460 20435 5500 20890
rect 5830 20445 5870 20970
rect 5920 20445 5960 21050
rect 6270 20445 6310 21130
rect 6475 20445 6515 21215
rect 6575 20445 6615 21305
rect 6940 20445 6980 21395
rect 7230 20445 7270 21485
rect 7325 20460 7365 21575
rect 7600 20435 7640 21665
rect 7710 20440 7750 21755
rect 7875 21715 7915 22385
rect 7870 21710 7920 21715
rect 7870 21670 7875 21710
rect 7915 21670 7920 21710
rect 7870 21665 7920 21670
rect 8025 21445 8065 22550
rect 8311 22495 8341 22576
rect 8020 21440 8070 21445
rect 8020 21400 8025 21440
rect 8065 21400 8070 21440
rect 8020 21395 8070 21400
rect 8305 21180 8345 22495
rect 8587 22490 8617 22576
rect 8863 22490 8893 22576
rect 9139 22490 9169 22576
rect 9415 22490 9445 22576
rect 8300 21175 8350 21180
rect 8300 21135 8305 21175
rect 8345 21135 8350 21175
rect 8300 21130 8350 21135
rect 8585 20940 8625 22490
rect 8860 22345 8900 22490
rect 8855 22340 8905 22345
rect 8855 22300 8860 22340
rect 8900 22300 8905 22340
rect 8855 22295 8905 22300
rect 9135 22075 9175 22490
rect 9130 22070 9180 22075
rect 9130 22030 9135 22070
rect 9175 22030 9180 22070
rect 9130 22025 9180 22030
rect 8580 20935 8630 20940
rect 8580 20895 8585 20935
rect 8625 20895 8630 20935
rect 8580 20890 8630 20895
rect 9410 20700 9450 22490
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22490 10273 22576
rect 10240 21625 10280 22490
rect 10519 22485 10549 22576
rect 10795 22490 10825 22576
rect 10235 21620 10285 21625
rect 10235 21580 10240 21620
rect 10280 21580 10285 21620
rect 10235 21575 10285 21580
rect 10515 21535 10555 22485
rect 10510 21530 10560 21535
rect 10510 21490 10515 21530
rect 10555 21490 10560 21530
rect 10510 21485 10560 21490
rect 10790 21355 10830 22490
rect 11071 22485 11101 22576
rect 11347 22490 11377 22576
rect 10785 21350 10835 21355
rect 10785 21310 10790 21350
rect 10830 21310 10835 21350
rect 10785 21305 10835 21310
rect 11065 21265 11105 22485
rect 11060 21260 11110 21265
rect 11060 21220 11065 21260
rect 11105 21220 11110 21260
rect 11060 21215 11110 21220
rect 11345 21100 11385 22490
rect 11623 22485 11653 22576
rect 11899 22490 11929 22576
rect 12175 22490 12205 22576
rect 12451 22490 12481 22576
rect 12727 22490 12757 22576
rect 11340 21095 11390 21100
rect 11340 21055 11345 21095
rect 11385 21055 11390 21095
rect 11340 21050 11390 21055
rect 11620 21020 11660 22485
rect 11615 21015 11665 21020
rect 11615 20975 11620 21015
rect 11660 20975 11665 21015
rect 11615 20970 11665 20975
rect 11895 20860 11935 22490
rect 11890 20855 11940 20860
rect 11890 20815 11895 20855
rect 11935 20815 11940 20855
rect 11890 20810 11940 20815
rect 12170 20780 12210 22490
rect 12445 22255 12485 22490
rect 12440 22250 12490 22255
rect 12440 22210 12445 22250
rect 12485 22210 12490 22250
rect 12440 22205 12490 22210
rect 12725 22165 12765 22490
rect 13003 22485 13033 22576
rect 13279 22485 13309 22576
rect 13555 22530 13585 22576
rect 12720 22160 12770 22165
rect 12720 22120 12725 22160
rect 12765 22120 12770 22160
rect 12720 22115 12770 22120
rect 13000 21985 13040 22485
rect 12995 21980 13045 21985
rect 12995 21940 13000 21980
rect 13040 21940 13045 21980
rect 12995 21935 13045 21940
rect 13275 21895 13315 22485
rect 13270 21890 13320 21895
rect 13270 21850 13275 21890
rect 13315 21850 13320 21890
rect 13270 21845 13320 21850
rect 12165 20775 12215 20780
rect 12165 20735 12170 20775
rect 12210 20735 12215 20775
rect 12165 20730 12215 20735
rect 9405 20695 9455 20700
rect 9405 20655 9410 20695
rect 9450 20655 9455 20695
rect 9405 20650 9455 20655
rect 13545 20620 13585 22530
rect 13831 22490 13861 22576
rect 13540 20615 13590 20620
rect 13540 20575 13545 20615
rect 13585 20575 13590 20615
rect 13540 20570 13590 20575
rect 13825 20540 13865 22490
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 13820 20535 13870 20540
rect 13820 20495 13825 20535
rect 13865 20495 13870 20535
rect 13820 20490 13870 20495
rect 400 19445 410 19485
rect 450 19445 475 19485
rect 515 19445 540 19485
rect 580 19445 600 19485
rect 400 500 600 19445
use add  add_0
timestamp 1747071801
transform 1 0 3080 0 1 20135
box -85 -695 4790 335
<< labels >>
flabel metal4 s 14383 22476 14413 22576 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 14659 22476 14689 22576 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 14107 22476 14137 22576 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 13831 22476 13861 22576 0 FreeSans 240 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 13555 22476 13585 22576 0 FreeSans 240 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 13279 22476 13309 22576 0 FreeSans 240 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 13003 22476 13033 22576 0 FreeSans 240 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 12727 22476 12757 22576 0 FreeSans 240 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 12451 22476 12481 22576 0 FreeSans 240 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 12175 22476 12205 22576 0 FreeSans 240 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 11899 22476 11929 22576 0 FreeSans 240 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 11623 22476 11653 22576 0 FreeSans 240 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 11347 22476 11377 22576 0 FreeSans 240 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 11071 22476 11101 22576 0 FreeSans 240 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 10795 22476 10825 22576 0 FreeSans 240 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 10519 22476 10549 22576 0 FreeSans 240 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 10243 22476 10273 22576 0 FreeSans 240 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 9967 22476 9997 22576 0 FreeSans 240 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 9691 22476 9721 22576 0 FreeSans 240 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 4999 22476 5029 22576 0 FreeSans 240 90 0 0 uio_oe[0]
port 19 nsew signal tristate
flabel metal4 s 4723 22476 4753 22576 0 FreeSans 240 90 0 0 uio_oe[1]
port 20 nsew signal tristate
flabel metal4 s 4447 22476 4477 22576 0 FreeSans 240 90 0 0 uio_oe[2]
port 21 nsew signal tristate
flabel metal4 s 4171 22476 4201 22576 0 FreeSans 240 90 0 0 uio_oe[3]
port 22 nsew signal tristate
flabel metal4 s 3895 22476 3925 22576 0 FreeSans 240 90 0 0 uio_oe[4]
port 23 nsew signal tristate
flabel metal4 s 3619 22476 3649 22576 0 FreeSans 240 90 0 0 uio_oe[5]
port 24 nsew signal tristate
flabel metal4 s 3343 22476 3373 22576 0 FreeSans 240 90 0 0 uio_oe[6]
port 25 nsew signal tristate
flabel metal4 s 3067 22476 3097 22576 0 FreeSans 240 90 0 0 uio_oe[7]
port 26 nsew signal tristate
flabel metal4 s 7207 22476 7237 22576 0 FreeSans 240 90 0 0 uio_out[0]
port 27 nsew signal tristate
flabel metal4 s 6931 22476 6961 22576 0 FreeSans 240 90 0 0 uio_out[1]
port 28 nsew signal tristate
flabel metal4 s 6655 22476 6685 22576 0 FreeSans 240 90 0 0 uio_out[2]
port 29 nsew signal tristate
flabel metal4 s 6379 22476 6409 22576 0 FreeSans 240 90 0 0 uio_out[3]
port 30 nsew signal tristate
flabel metal4 s 6103 22476 6133 22576 0 FreeSans 240 90 0 0 uio_out[4]
port 31 nsew signal tristate
flabel metal4 s 5827 22476 5857 22576 0 FreeSans 240 90 0 0 uio_out[5]
port 32 nsew signal tristate
flabel metal4 s 5551 22476 5581 22576 0 FreeSans 240 90 0 0 uio_out[6]
port 33 nsew signal tristate
flabel metal4 s 5275 22476 5305 22576 0 FreeSans 240 90 0 0 uio_out[7]
port 34 nsew signal tristate
flabel metal4 s 9415 22476 9445 22576 0 FreeSans 240 90 0 0 uo_out[0]
port 35 nsew signal tristate
flabel metal4 s 9139 22476 9169 22576 0 FreeSans 240 90 0 0 uo_out[1]
port 36 nsew signal tristate
flabel metal4 s 8863 22476 8893 22576 0 FreeSans 240 90 0 0 uo_out[2]
port 37 nsew signal tristate
flabel metal4 s 8587 22476 8617 22576 0 FreeSans 240 90 0 0 uo_out[3]
port 38 nsew signal tristate
flabel metal4 s 8311 22476 8341 22576 0 FreeSans 240 90 0 0 uo_out[4]
port 39 nsew signal tristate
flabel metal4 s 8035 22476 8065 22576 0 FreeSans 240 90 0 0 uo_out[5]
port 40 nsew signal tristate
flabel metal4 s 7759 22476 7789 22576 0 FreeSans 240 90 0 0 uo_out[6]
port 41 nsew signal tristate
flabel metal4 s 7483 22476 7513 22576 0 FreeSans 240 90 0 0 uo_out[7]
port 42 nsew signal tristate
flabel metal4 100 500 300 22076 1 FreeSans 1 0 0 0 VDPWR
port 43 nsew power bidirectional
flabel metal4 400 500 600 22076 1 FreeSans 1 0 0 0 VGND
port 44 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
