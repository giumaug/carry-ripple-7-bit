VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO test
  CLASS BLOCK ;
  FOREIGN test ;
  ORIGIN -1.000 -5.000 ;
  SIZE 293.000 BY 220.760 ;
  OBS
      LAYER met3 ;
        RECT 1.000 187.000 294.000 220.000 ;
      LAYER met4 ;
        RECT 1.000 5.000 277.300 225.760 ;
  END
END test
END LIBRARY

