* NGSPICE file created from tt_um_carry_ripple_7_bit.ext - technology: sky130A

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.177 ps=1.69 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.138 ps=1.4 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.69 as=0.177 ps=1.69 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.4 as=0.0878 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.4 as=0.25 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.69 as=0.177 ps=1.69 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.69 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.138 ps=1.4 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.103 pd=0.954 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.245 ps=2.27 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.816 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.103 ps=0.954 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.136 ps=1.26 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.229 ps=1.57 w=0.65 l=0.15
**devattr s=10270,288 d=3575,185
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5500,255
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.18 ps=1.69 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.229 pd=1.57 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=10270,288
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.229 pd=1.57 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=6890,366
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.18 ps=1.69 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
**devattr s=3575,185 d=3640,186
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.226 ps=2.26 w=0.87 l=1.97
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=1.97
**devattr d=5720,324
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.226 pd=2.26 as=0.226 ps=2.26 w=0.87 l=1.05
**devattr d=9048,452
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.143 ps=1.62 w=0.55 l=1.05
**devattr d=5720,324
.ends

.subckt add A1 B1 CI S1 A2 B2 S2 A3 B3 S3 A4 B4 S4 A5 B5 S5 A6 B6 S6 A7 B7 S7 CO VDD_1
+ VDD_2 VDD_3 sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__xor2_1_9/VPB VSUBS
Xsky130_fd_sc_hd__xor2_1_3 A4 B4 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__xor2_1_3/X sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_4 A5 B5 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__xor2_1_4/X sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_5 A6 sky130_fd_sc_hd__xor2_1_5/B VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__xor2_1_5/X sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_6 A7 B7 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__xor2_1_6/X sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_7 sky130_fd_sc_hd__xor2_1_7/A CI VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB
+ sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_7/X sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_8 sky130_fd_sc_hd__xor2_1_8/A sky130_fd_sc_hd__xor2_1_8/B
+ VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_8/X
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_1_0 A1 sky130_fd_sc_hd__and2_1_0/B VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__and2_1_0/X sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__xor2_1_9 sky130_fd_sc_hd__xor2_1_9/A sky130_fd_sc_hd__xor2_1_9/B
+ VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/X
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_1_1 A2 sky130_fd_sc_hd__and2_1_1/B VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__and2_1_1/X sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_3 A4 B4 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__and2_1_3/X sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_2 A3 B3 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__and2_1_2/X sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_4 A5 B5 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__and2_1_4/X sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_5 A6 sky130_fd_sc_hd__xor2_1_5/B VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__and2_1_5/X sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_6 A7 B7 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__and2_1_6/X sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__a21o_1_0 sky130_fd_sc_hd__xor2_1_7/A sky130_fd_sc_hd__a21o_1_0/A2
+ sky130_fd_sc_hd__and2_1_0/X VSUBS VSUBS VDD_2 VDD_2 sky130_fd_sc_hd__a21o_1_0/X
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_2 sky130_fd_sc_hd__xor2_1_9/A sky130_fd_sc_hd__xor2_1_9/B
+ sky130_fd_sc_hd__and2_1_2/X VSUBS VSUBS VDD_2 VDD_2 sky130_fd_sc_hd__a21o_1_2/X
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_1 sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__xor2_1_1/X
+ sky130_fd_sc_hd__and2_1_1/X VSUBS VSUBS VDD_2 VDD_2 sky130_fd_sc_hd__xor2_1_9/A
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_3 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__xor2_1_3/X
+ sky130_fd_sc_hd__and2_1_3/X VSUBS VSUBS VDD_2 VDD_2 sky130_fd_sc_hd__a21o_1_3/X
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_4 sky130_fd_sc_hd__a21o_1_3/X sky130_fd_sc_hd__xor2_1_4/X
+ sky130_fd_sc_hd__a21o_1_4/B1 VSUBS VSUBS VDD_2 VDD_2 sky130_fd_sc_hd__a21o_1_4/X
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_5 sky130_fd_sc_hd__xor2_1_12/A sky130_fd_sc_hd__xor2_1_5/X
+ sky130_fd_sc_hd__and2_1_5/X VSUBS VSUBS VDD_2 VDD_2 sky130_fd_sc_hd__a21o_1_5/X
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_6 sky130_fd_sc_hd__a21o_1_5/X sky130_fd_sc_hd__xor2_1_6/X
+ sky130_fd_sc_hd__and2_1_6/X VSUBS VSUBS VDD_2 VDD_2 CO sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__decap_6_0 VSUBS VSUBS VDD_2 VDD_2 sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_1 VSUBS VSUBS VDD_2 VDD_2 sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_2 VSUBS VSUBS VDD_2 VDD_2 sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_3 VSUBS VSUBS VDD_2 VDD_2 sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_4_0 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/VPB
+ sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_6_5 VSUBS VSUBS VDD_2 VDD_2 sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_4 VSUBS VSUBS VDD_2 VDD_2 sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_4_1 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/VPB
+ sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_6_6 VSUBS VSUBS VDD_2 VDD_2 sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_4_2 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/VPB
+ sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__xor2_1_10 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__xor2_1_3/X
+ VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/VPB S4 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_6_7 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/VPB
+ sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__xor2_1_11 sky130_fd_sc_hd__xor2_1_4/X sky130_fd_sc_hd__a21o_1_3/X
+ VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/VPB S5 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_6_8 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/VPB
+ sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__xor2_1_12 sky130_fd_sc_hd__xor2_1_12/A sky130_fd_sc_hd__xor2_1_5/X
+ VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/VPB S6 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_6_9 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/VPB
+ sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__xor2_1_13 sky130_fd_sc_hd__xor2_1_6/X sky130_fd_sc_hd__a21o_1_5/X
+ VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/VPB S7 sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__decap_6_10 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_9/VPB sky130_fd_sc_hd__xor2_1_9/VPB
+ sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__xor2_1_0 A1 sky130_fd_sc_hd__xor2_1_0/B VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_2 A3 sky130_fd_sc_hd__xor2_1_2/B VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__xor2_1_2/X sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_1 A2 B2 VSUBS VSUBS sky130_fd_sc_hd__xor2_1_6/VPB sky130_fd_sc_hd__xor2_1_6/VPB
+ sky130_fd_sc_hd__xor2_1_1/X sky130_fd_sc_hd__xor2_1
.ends

.subckt tt_um_carry_ripple_7_bit clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] VDPWR VGND
Xadd_0 ui_in[0] ui_in[1] VGND uo_out[0] ui_in[2] ui_in[3] uo_out[1] ui_in[4] ui_in[5]
+ uo_out[2] ui_in[6] ui_in[7] uo_out[3] uio_in[0] uio_in[1] uo_out[4] uio_in[2] uio_in[3]
+ uo_out[5] uio_in[4] uio_in[5] uo_out[6] uo_out[7] VDPWR VDPWR VDPWR VDPWR VDPWR
+ VGND add
.ends

