magic
tech sky130A
magscale 1 2
timestamp 1738491202
<< metal1 >>
rect 1816 18235 6940 18350
rect 7260 18190 7350 18200
rect 7260 18120 7270 18190
rect 7340 18120 7350 18190
rect 8540 18190 8630 18200
rect 9980 18190 10070 18200
rect 8540 18120 8550 18190
rect 8620 18120 8630 18190
rect 7260 18110 7350 18120
rect 8020 18110 8110 18120
rect 8540 18110 8630 18120
rect 9290 18180 9390 18190
rect 9290 18110 9300 18180
rect 9380 18110 9390 18180
rect 9980 18120 9990 18190
rect 10060 18120 10070 18190
rect 11260 18190 11350 18200
rect 11260 18120 11270 18190
rect 11340 18120 11350 18190
rect 9980 18110 10070 18120
rect 10730 18110 10820 18120
rect 11260 18110 11350 18120
rect 12010 18170 12100 18180
rect 7030 18030 7050 18070
rect 8020 18040 8030 18110
rect 8100 18040 8110 18110
rect 9290 18100 9390 18110
rect 8020 18030 8110 18040
rect 10730 18040 10740 18110
rect 10810 18040 10820 18110
rect 12010 18100 12020 18170
rect 12090 18100 12100 18170
rect 12010 18090 12100 18100
rect 10730 18030 10820 18040
rect 6960 18020 7050 18030
rect 10490 18020 10580 18030
rect 6960 17950 6970 18020
rect 7040 17950 7050 18020
rect 6960 17940 7050 17950
rect 7530 18010 7620 18020
rect 7530 17940 7540 18010
rect 7610 17940 7620 18010
rect 7530 17930 7620 17940
rect 8240 18010 8330 18020
rect 8240 17940 8250 18010
rect 8320 17940 8330 18010
rect 8240 17930 8330 17940
rect 8810 18010 8900 18020
rect 8810 17940 8820 18010
rect 8890 17940 8900 18010
rect 8810 17930 8900 17940
rect 9680 18010 9770 18020
rect 9680 17940 9690 18010
rect 9680 17930 9770 17940
rect 10490 17950 10500 18020
rect 10570 17950 10580 18020
rect 10490 17940 10580 17950
rect 10960 18010 11050 18020
rect 10960 17940 10970 18010
rect 11040 17940 11050 18010
rect 8810 17900 8830 17930
rect 8890 17890 8900 17930
rect 10490 17900 10510 17940
rect 10960 17930 11050 17940
rect 11520 18000 11610 18020
rect 11520 17930 11530 18000
rect 11600 17930 11610 18000
rect 11520 17900 11550 17930
rect 11590 17890 11610 17930
rect 1816 17690 6935 17805
<< via1 >>
rect 7270 18120 7340 18190
rect 8550 18120 8620 18190
rect 9300 18110 9380 18180
rect 9990 18120 10060 18190
rect 11270 18120 11340 18190
rect 8030 18040 8100 18110
rect 10740 18040 10810 18110
rect 12020 18100 12090 18170
rect 6970 17950 7040 18020
rect 7540 17940 7610 18010
rect 8250 17940 8320 18010
rect 8820 17940 8890 18010
rect 9690 17940 9770 18010
rect 10500 17950 10570 18020
rect 10970 17940 11040 18010
rect 11530 17930 11600 18000
<< metal2 >>
rect 11520 21650 11610 21660
rect 11520 21570 11530 21650
rect 11600 21570 11610 21650
rect 11520 21560 11610 21570
rect 10950 21470 11040 21480
rect 10950 21390 10960 21470
rect 11030 21390 11040 21470
rect 10950 21380 11040 21390
rect 10500 21290 10580 21300
rect 10500 21230 10510 21290
rect 10570 21230 10580 21290
rect 10500 21220 10580 21230
rect 9680 21120 9770 21140
rect 9680 21050 9700 21120
rect 9760 21050 9770 21120
rect 9680 21040 9770 21050
rect 8810 20940 8890 20960
rect 8810 20880 8820 20940
rect 8880 20880 8890 20940
rect 8810 20860 8890 20880
rect 8260 20760 8340 20780
rect 8260 20690 8270 20760
rect 8330 20690 8340 20760
rect 8260 20680 8340 20690
rect 7540 20580 7620 20600
rect 7540 20520 7550 20580
rect 7610 20520 7620 20580
rect 7540 20500 7620 20520
rect 6970 20400 7050 20420
rect 6970 20340 6980 20400
rect 7040 20340 7050 20400
rect 6970 20320 7050 20340
rect 6980 18030 7030 20320
rect 7260 18960 7340 18980
rect 7260 18900 7270 18960
rect 7330 18900 7340 18960
rect 7260 18880 7340 18900
rect 7270 18200 7320 18880
rect 7260 18190 7350 18200
rect 7260 18120 7270 18190
rect 7340 18120 7350 18190
rect 7260 18110 7350 18120
rect 6960 18020 7050 18030
rect 7550 18020 7600 20500
rect 8020 19140 8100 19160
rect 8020 19080 8030 19140
rect 8090 19080 8100 19140
rect 8020 19060 8100 19080
rect 8030 18120 8080 19060
rect 8020 18110 8110 18120
rect 8020 18040 8030 18110
rect 8100 18040 8110 18110
rect 8020 18030 8110 18040
rect 8270 18020 8320 20680
rect 8550 19320 8630 19340
rect 8550 19260 8560 19320
rect 8620 19260 8630 19320
rect 8550 19240 8630 19260
rect 8560 18200 8610 19240
rect 8540 18190 8630 18200
rect 8540 18120 8550 18190
rect 8620 18120 8630 18190
rect 8540 18110 8630 18120
rect 8830 18020 8880 20860
rect 9300 19500 9380 19520
rect 9300 19440 9310 19500
rect 9370 19440 9380 19500
rect 9300 19420 9380 19440
rect 9310 18190 9360 19420
rect 9290 18180 9390 18190
rect 9290 18110 9300 18180
rect 9380 18110 9390 18180
rect 9290 18100 9390 18110
rect 9700 18020 9760 21040
rect 9990 19680 10070 19700
rect 9990 19620 10000 19680
rect 10060 19620 10070 19680
rect 9990 19600 10070 19620
rect 10000 18200 10050 19600
rect 9980 18190 10070 18200
rect 9980 18120 9990 18190
rect 10060 18120 10070 18190
rect 9980 18110 10070 18120
rect 10520 18030 10570 21220
rect 10970 20240 11030 21380
rect 10740 19860 10820 19880
rect 10740 19800 10750 19860
rect 10810 19800 10820 19860
rect 10740 19780 10820 19800
rect 10750 18120 10800 19780
rect 10972 18578 11030 20240
rect 11270 20040 11350 20060
rect 11270 19980 11280 20040
rect 11340 19980 11350 20040
rect 11270 19960 11350 19980
rect 10970 18348 11030 18578
rect 10730 18110 10820 18120
rect 10730 18040 10740 18110
rect 10810 18040 10820 18110
rect 10730 18030 10820 18040
rect 10490 18020 10580 18030
rect 10978 18020 11028 18348
rect 11280 18200 11330 19960
rect 11260 18190 11350 18200
rect 11260 18120 11270 18190
rect 11340 18120 11350 18190
rect 11260 18110 11350 18120
rect 6960 17950 6970 18020
rect 7040 17950 7050 18020
rect 6960 17940 7050 17950
rect 7530 18010 7620 18020
rect 7530 17940 7540 18010
rect 7610 17940 7620 18010
rect 7530 17930 7620 17940
rect 8240 18010 8330 18020
rect 8240 17940 8250 18010
rect 8320 17940 8330 18010
rect 8240 17930 8330 17940
rect 8810 18010 8900 18020
rect 8810 17940 8820 18010
rect 8890 17940 8900 18010
rect 8810 17930 8900 17940
rect 9680 18010 9780 18020
rect 9680 17940 9690 18010
rect 9770 17940 9780 18010
rect 10490 17950 10500 18020
rect 10570 17950 10580 18020
rect 10490 17940 10580 17950
rect 10960 18010 11050 18020
rect 11540 18010 11590 21560
rect 12020 20220 12100 20240
rect 12020 20160 12030 20220
rect 12090 20160 12100 20220
rect 12020 20140 12100 20160
rect 12030 18180 12080 20140
rect 12010 18170 12100 18180
rect 12010 18100 12020 18170
rect 12090 18100 12100 18170
rect 12010 18090 12100 18100
rect 10960 17940 10970 18010
rect 11040 17940 11050 18010
rect 9680 17930 9780 17940
rect 10960 17930 11050 17940
rect 11520 18000 11610 18010
rect 11520 17930 11530 18000
rect 11600 17930 11610 18000
rect 11520 17920 11610 17930
<< via2 >>
rect 11530 21570 11600 21650
rect 10960 21390 11030 21470
rect 10510 21230 10570 21290
rect 9700 21050 9760 21120
rect 8820 20880 8880 20940
rect 8270 20690 8330 20760
rect 7550 20520 7610 20580
rect 6980 20340 7040 20400
rect 7270 18900 7330 18960
rect 8030 19080 8090 19140
rect 8560 19260 8620 19320
rect 9310 19440 9370 19500
rect 10000 19620 10060 19680
rect 10750 19800 10810 19860
rect 11280 19980 11340 20040
rect 12030 20160 12090 20220
<< metal3 >>
rect 1816 21830 29400 21840
rect 1816 21750 6130 21830
rect 6200 21750 6680 21830
rect 6750 21750 7230 21830
rect 7300 21750 7780 21830
rect 7850 21750 8340 21830
rect 8410 21750 8890 21830
rect 8960 21750 9440 21830
rect 9510 21750 9990 21830
rect 10060 21750 10540 21830
rect 10610 21750 11100 21830
rect 11170 21750 11650 21830
rect 11720 21750 12200 21830
rect 12270 21750 12750 21830
rect 12820 21750 13300 21830
rect 13370 21750 13860 21830
rect 13930 21750 14410 21830
rect 14480 21750 29400 21830
rect 1816 21740 29400 21750
rect 6080 21650 29400 21660
rect 6080 21570 11530 21650
rect 11600 21570 23780 21650
rect 23860 21570 29400 21650
rect 6080 21560 29400 21570
rect 6080 21470 29400 21480
rect 6080 21390 10960 21470
rect 11030 21390 24340 21470
rect 24410 21390 29400 21470
rect 6080 21380 29400 21390
rect 24880 21300 24990 21310
rect 6080 21290 24880 21300
rect 6080 21230 10510 21290
rect 10570 21230 24880 21290
rect 6080 21220 24880 21230
rect 24980 21220 29400 21300
rect 24880 21210 24990 21220
rect 6080 21130 29400 21140
rect 6080 21120 25450 21130
rect 6080 21050 9700 21120
rect 9760 21050 25450 21120
rect 6080 21048 25450 21050
rect 25530 21048 29400 21130
rect 6080 21040 29400 21048
rect 6080 20950 29400 20960
rect 6080 20940 26000 20950
rect 6080 20880 8820 20940
rect 8880 20880 26000 20940
rect 6080 20870 26000 20880
rect 26080 20870 29400 20950
rect 6080 20860 29400 20870
rect 6080 20770 29400 20780
rect 6080 20760 26540 20770
rect 6080 20690 8270 20760
rect 8330 20690 26540 20760
rect 26620 20690 29400 20770
rect 6080 20680 29400 20690
rect 6080 20590 29400 20600
rect 6080 20580 27100 20590
rect 6080 20520 7550 20580
rect 7610 20520 27100 20580
rect 6080 20510 27100 20520
rect 27180 20510 29400 20590
rect 6080 20500 29400 20510
rect 6080 20410 29400 20420
rect 6080 20400 27640 20410
rect 6080 20340 6980 20400
rect 7040 20340 27640 20400
rect 6080 20330 27640 20340
rect 27720 20330 29400 20410
rect 6080 20320 29400 20330
rect 6080 20230 29400 20240
rect 6080 20220 14960 20230
rect 6080 20160 12030 20220
rect 12090 20160 14960 20220
rect 6080 20150 14960 20160
rect 15030 20150 29400 20230
rect 6080 20140 29400 20150
rect 6080 20050 29400 20060
rect 6080 20040 15510 20050
rect 6080 19980 11280 20040
rect 11340 19980 15510 20040
rect 6080 19970 15510 19980
rect 15580 19970 29400 20050
rect 6080 19960 29400 19970
rect 6080 19870 29400 19880
rect 6080 19860 16060 19870
rect 6080 19800 10750 19860
rect 10810 19800 16060 19860
rect 6080 19790 16060 19800
rect 16130 19790 29400 19870
rect 6080 19780 29400 19790
rect 6080 19690 29400 19700
rect 6080 19680 16620 19690
rect 6080 19620 10000 19680
rect 10060 19620 16620 19680
rect 6080 19610 16620 19620
rect 16690 19610 29400 19690
rect 6080 19600 29400 19610
rect 6080 19510 29400 19520
rect 6080 19500 17160 19510
rect 6080 19440 9310 19500
rect 9370 19440 17160 19500
rect 6080 19430 17160 19440
rect 17240 19430 29400 19510
rect 6080 19420 29400 19430
rect 6080 19330 29400 19340
rect 6080 19320 17720 19330
rect 6080 19260 8560 19320
rect 8620 19260 17720 19320
rect 6080 19250 17720 19260
rect 17800 19250 29400 19330
rect 6080 19240 29400 19250
rect 6080 19150 29400 19160
rect 6080 19140 18260 19150
rect 6080 19080 8030 19140
rect 8090 19080 18260 19140
rect 6080 19070 18260 19080
rect 18340 19070 29400 19150
rect 6080 19060 29400 19070
rect 6080 18970 29400 18980
rect 6080 18960 18820 18970
rect 6080 18900 7270 18960
rect 7330 18900 18820 18960
rect 6080 18890 18820 18900
rect 18900 18890 29400 18970
rect 6080 18880 29400 18890
rect 6080 18700 29400 18800
<< via3 >>
rect 6130 21750 6200 21830
rect 6680 21750 6750 21830
rect 7230 21750 7300 21830
rect 7780 21750 7850 21830
rect 8340 21750 8410 21830
rect 8890 21750 8960 21830
rect 9440 21750 9510 21830
rect 9990 21750 10060 21830
rect 10540 21750 10610 21830
rect 11100 21750 11170 21830
rect 11650 21750 11720 21830
rect 12200 21750 12270 21830
rect 12750 21750 12820 21830
rect 13300 21750 13370 21830
rect 13860 21750 13930 21830
rect 14410 21750 14480 21830
rect 23780 21570 23860 21650
rect 24340 21390 24410 21470
rect 24880 21220 24980 21300
rect 25450 21048 25530 21130
rect 26000 20870 26080 20950
rect 26540 20690 26620 20770
rect 27100 20510 27180 20590
rect 27640 20330 27720 20410
rect 14960 20150 15030 20230
rect 15510 19970 15580 20050
rect 16060 19790 16130 19870
rect 16620 19610 16690 19690
rect 17160 19430 17240 19510
rect 17720 19250 17800 19330
rect 18260 19070 18340 19150
rect 18820 18890 18900 18970
<< metal4 >>
rect 6120 21840 6200 21928
rect 6680 21840 6750 21928
rect 7230 21840 7300 21928
rect 7780 21840 7850 21928
rect 8340 21840 8410 21928
rect 8890 21840 8960 21928
rect 9440 21840 9510 21928
rect 9990 21840 10060 21928
rect 10540 21840 10610 21928
rect 11100 21840 11170 21928
rect 11650 21840 11720 21928
rect 12200 21840 12270 21928
rect 12750 21840 12820 21934
rect 13300 21840 13370 21934
rect 13860 21840 13930 21934
rect 14410 21840 14480 21934
rect 6110 21830 6210 21840
rect 6110 21750 6130 21830
rect 6200 21750 6210 21830
rect 6110 21740 6210 21750
rect 6660 21830 6760 21840
rect 6660 21750 6680 21830
rect 6750 21750 6760 21830
rect 6660 21740 6760 21750
rect 7210 21830 7310 21840
rect 7210 21750 7230 21830
rect 7300 21750 7310 21830
rect 7210 21740 7310 21750
rect 7760 21830 7860 21840
rect 7760 21750 7780 21830
rect 7850 21750 7860 21830
rect 7760 21740 7860 21750
rect 8320 21830 8420 21840
rect 8320 21750 8340 21830
rect 8410 21750 8420 21830
rect 8320 21740 8420 21750
rect 8870 21830 8970 21840
rect 8870 21750 8890 21830
rect 8960 21750 8970 21830
rect 8870 21740 8970 21750
rect 9420 21830 9520 21840
rect 9420 21750 9440 21830
rect 9510 21750 9520 21830
rect 9420 21740 9520 21750
rect 9970 21830 10070 21840
rect 9970 21750 9990 21830
rect 10060 21750 10070 21830
rect 9970 21740 10070 21750
rect 10520 21830 10620 21840
rect 10520 21750 10540 21830
rect 10610 21750 10620 21830
rect 10520 21740 10620 21750
rect 11080 21830 11180 21840
rect 11080 21750 11100 21830
rect 11170 21750 11180 21830
rect 11080 21740 11180 21750
rect 11630 21830 11730 21840
rect 11630 21750 11650 21830
rect 11720 21750 11730 21830
rect 11630 21740 11730 21750
rect 12180 21830 12280 21840
rect 12180 21750 12200 21830
rect 12270 21750 12280 21830
rect 12180 21740 12280 21750
rect 12730 21830 12830 21840
rect 12730 21750 12750 21830
rect 12820 21750 12830 21830
rect 12730 21740 12830 21750
rect 13280 21830 13380 21840
rect 13280 21750 13300 21830
rect 13370 21750 13380 21830
rect 13280 21740 13380 21750
rect 13840 21830 13940 21840
rect 13840 21750 13860 21830
rect 13930 21750 13940 21830
rect 13840 21740 13940 21750
rect 14390 21830 14490 21840
rect 14390 21750 14410 21830
rect 14480 21750 14490 21830
rect 14390 21740 14490 21750
rect 14960 20240 15030 21934
rect 14950 20230 15040 20240
rect 14950 20150 14960 20230
rect 15030 20150 15040 20230
rect 14950 20140 15040 20150
rect 15510 20060 15580 21934
rect 15500 20050 15590 20060
rect 15500 19970 15510 20050
rect 15580 19970 15590 20050
rect 15500 19960 15590 19970
rect 16060 19880 16130 21934
rect 16050 19870 16140 19880
rect 16050 19790 16060 19870
rect 16130 19790 16140 19870
rect 16050 19780 16140 19790
rect 16620 19700 16690 21934
rect 16610 19690 16700 19700
rect 16610 19610 16620 19690
rect 16690 19610 16700 19690
rect 16610 19600 16700 19610
rect 17160 19520 17240 21934
rect 17150 19510 17250 19520
rect 17150 19430 17160 19510
rect 17240 19430 17250 19510
rect 17150 19420 17250 19430
rect 17720 19340 17800 21934
rect 17710 19330 17810 19340
rect 17710 19250 17720 19330
rect 17800 19250 17810 19330
rect 17710 19240 17810 19250
rect 18260 19160 18340 21934
rect 18250 19150 18350 19160
rect 18250 19070 18260 19150
rect 18340 19070 18350 19150
rect 18250 19060 18350 19070
rect 18820 18980 18900 21934
rect 23790 21660 23860 21934
rect 23770 21650 23870 21660
rect 23770 21570 23780 21650
rect 23860 21570 23870 21650
rect 23770 21560 23870 21570
rect 24350 21480 24410 21934
rect 24330 21470 24420 21480
rect 24330 21390 24340 21470
rect 24410 21390 24420 21470
rect 24330 21380 24420 21390
rect 24900 21310 24970 21934
rect 24870 21300 24990 21310
rect 24870 21220 24880 21300
rect 24980 21220 24990 21300
rect 24870 21210 24990 21220
rect 25450 21140 25530 21934
rect 25430 21130 25540 21140
rect 25430 21048 25450 21130
rect 25530 21048 25540 21130
rect 25430 21040 25540 21048
rect 26000 20960 26080 21934
rect 25980 20950 26090 20960
rect 25980 20870 26000 20950
rect 26080 20870 26090 20950
rect 25980 20860 26090 20870
rect 26540 20780 26620 21934
rect 26520 20770 26630 20780
rect 26520 20690 26540 20770
rect 26620 20690 26630 20770
rect 26520 20680 26630 20690
rect 27100 20600 27180 21934
rect 27080 20590 27190 20600
rect 27080 20510 27100 20590
rect 27180 20510 27190 20590
rect 27080 20500 27190 20510
rect 27640 20420 27720 21934
rect 27620 20410 27730 20420
rect 27620 20330 27640 20410
rect 27720 20330 27730 20410
rect 27620 20320 27730 20330
rect 18810 18970 18910 18980
rect 18810 18890 18820 18970
rect 18900 18890 18910 18970
rect 18810 18880 18910 18890
use adder_1  adder_1_0
timestamp 1700079872
transform 1 0 6960 0 1 17750
box -80 -50 5188 590
<< labels >>
rlabel via3 6160 21768 6170 21806 1 PP1
port 1 n
rlabel via3 6694 21762 6728 21800 1 PP2
port 2 n
rlabel via3 7252 21766 7274 21800 1 PP3
port 3 n
rlabel via3 7790 21764 7810 21792 1 PP4
port 4 n
rlabel via3 8362 21780 8382 21808 1 PP5
port 5 n
rlabel via3 8908 21758 8932 21796 1 PP6
port 6 n
rlabel via3 9458 21776 9486 21808 1 PP7
port 7 n
rlabel via3 10024 21780 10052 21812 1 PP8
port 8 n
rlabel via3 10556 21788 10584 21820 1 PP9
port 9 n
rlabel via3 11110 21762 11134 21802 1 PP10
port 10 n
rlabel via3 11674 21788 11698 21828 1 PP11
port 11 n
rlabel via3 12208 21778 12228 21808 1 PP12
port 12 n
rlabel via3 12776 21796 12796 21826 1 PP13
port 13 n
rlabel via3 13330 21774 13350 21804 1 PP14
port 14 n
rlabel via3 13882 21792 13902 21822 1 PP15
port 15 n
rlabel via3 14438 21794 14458 21824 1 PP16
port 16 n
rlabel metal4 14970 21794 14990 21824 1 PP17
port 17 n
rlabel metal4 15524 21804 15544 21834 1 PP18
port 18 n
rlabel metal4 16084 21786 16104 21816 1 PP19
port 19 n
rlabel metal4 16640 21810 16660 21840 1 PP20
port 20 n
rlabel metal4 17194 21790 17214 21820 1 PP21
port 21 n
rlabel metal4 17746 21794 17766 21824 1 PP22
port 22 n
rlabel metal4 18294 21800 18314 21830 1 PP23
port 23 n
rlabel metal4 18840 21774 18860 21804 1 PP24
port 24 n
rlabel metal4 23818 21792 23838 21822 1 PP25
port 25 n
rlabel metal4 24384 21800 24404 21830 1 PP26
port 26 n
rlabel metal4 24922 21782 24942 21812 1 PP27
port 27 n
rlabel metal4 25474 21788 25494 21818 1 PP28
port 28 n
rlabel metal4 26022 21782 26042 21812 1 PP29
port 29 n
rlabel metal4 26576 21808 26596 21838 1 PP30
port 30 n
rlabel metal4 27152 21802 27172 21832 1 PP31
port 31 n
rlabel metal4 27670 21800 27690 21830 1 PP32
port 32 n
rlabel metal3 1958 21774 2016 21796 1 PP33
port 33 n
rlabel metal1 1844 18294 1902 18316 1 PP34
port 34 n
rlabel metal1 1920 17748 1978 17770 1 PP35
port 35 n
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
