magic
tech sky130A
magscale 1 2
timestamp 1738578133
<< metal3 >>
rect 400 21990 945 22000
rect 400 21950 410 21990
rect 450 21950 470 21990
rect 510 21950 530 21990
rect 570 21951 945 21990
rect 570 21950 600 21951
rect 815 21950 945 21951
rect 400 21935 600 21950
rect 100 20245 300 20255
rect 100 20205 110 20245
rect 150 20205 170 20245
rect 210 20205 230 20245
rect 270 20205 300 20245
rect 100 20195 300 20205
rect 400 19975 600 19985
rect 400 19935 410 19975
rect 450 19935 470 19975
rect 510 19935 530 19975
rect 570 19935 600 19975
rect 400 19925 600 19935
rect 1816 21830 29400 21840
rect 1816 21750 6130 21830
rect 6200 21750 6680 21830
rect 6750 21750 7230 21830
rect 7300 21750 7780 21830
rect 7850 21750 8340 21830
rect 8410 21750 8890 21830
rect 8960 21750 9440 21830
rect 9510 21750 9990 21830
rect 10060 21750 10540 21830
rect 10610 21750 11100 21830
rect 11170 21750 11650 21830
rect 11720 21750 12200 21830
rect 12270 21750 12750 21830
rect 12820 21750 13300 21830
rect 13370 21750 13860 21830
rect 13930 21750 14410 21830
rect 14480 21750 29400 21830
rect 1816 21740 29400 21750
rect 6080 21650 29400 21660
rect 6080 21570 11530 21650
rect 11600 21570 23780 21650
rect 23860 21570 29400 21650
rect 6080 21560 29400 21570
rect 6080 21470 29400 21480
rect 6080 21390 10960 21470
rect 11030 21390 24340 21470
rect 24410 21390 29400 21470
rect 6080 21380 29400 21390
rect 24880 21300 24990 21310
rect 6080 21290 24880 21300
rect 6080 21230 10510 21290
rect 10570 21230 24880 21290
rect 6080 21220 24880 21230
rect 24980 21220 29400 21300
rect 24880 21210 24990 21220
rect 6080 21130 29400 21140
rect 6080 21120 25450 21130
rect 6080 21050 9700 21120
rect 9760 21050 25450 21120
rect 6080 21048 25450 21050
rect 25530 21048 29400 21130
rect 6080 21040 29400 21048
rect 6080 20950 29400 20960
rect 6080 20940 26000 20950
rect 6080 20880 8820 20940
rect 8880 20880 26000 20940
rect 6080 20870 26000 20880
rect 26080 20870 29400 20950
rect 6080 20860 29400 20870
rect 6080 20770 29400 20780
rect 6080 20760 26540 20770
rect 6080 20690 8270 20760
rect 8330 20690 26540 20760
rect 26620 20690 29400 20770
rect 6080 20680 29400 20690
rect 6080 20590 29400 20600
rect 6080 20580 27100 20590
rect 6080 20520 7550 20580
rect 7610 20520 27100 20580
rect 6080 20510 27100 20520
rect 27180 20510 29400 20590
rect 6080 20500 29400 20510
rect 6080 20410 29400 20420
rect 6080 20400 27640 20410
rect 6080 20340 6980 20400
rect 7040 20340 27640 20400
rect 6080 20330 27640 20340
rect 27720 20330 29400 20410
rect 6080 20320 29400 20330
rect 6080 20230 29400 20240
rect 6080 20220 14960 20230
rect 6080 20160 12030 20220
rect 12090 20160 14960 20220
rect 6080 20150 14960 20160
rect 15030 20150 29400 20230
rect 6080 20140 29400 20150
rect 6080 20050 29400 20060
rect 6080 20040 15510 20050
rect 6080 19980 11280 20040
rect 11340 19980 15510 20040
rect 6080 19970 15510 19980
rect 15580 19970 29400 20050
rect 6080 19960 29400 19970
rect 6080 19870 29400 19880
rect 6080 19860 16060 19870
rect 6080 19800 10750 19860
rect 10810 19800 16060 19860
rect 6080 19790 16060 19800
rect 16130 19790 29400 19870
rect 6080 19780 29400 19790
rect 6080 19690 29400 19700
rect 6080 19680 16620 19690
rect 6080 19620 10000 19680
rect 10060 19620 16620 19680
rect 6080 19610 16620 19620
rect 16690 19610 29400 19690
rect 6080 19600 29400 19610
rect 6080 19510 29400 19520
rect 6080 19500 17160 19510
rect 6080 19440 9310 19500
rect 9370 19440 17160 19500
rect 6080 19430 17160 19440
rect 17240 19430 29400 19510
rect 6080 19420 29400 19430
rect 6080 19330 29400 19340
rect 6080 19320 17720 19330
rect 6080 19260 8560 19320
rect 8620 19260 17720 19320
rect 6080 19250 17720 19260
rect 17800 19250 29400 19330
rect 6080 19240 29400 19250
rect 6080 19150 29400 19160
rect 6080 19140 18260 19150
rect 6080 19080 8030 19140
rect 8090 19080 18260 19140
rect 6080 19070 18260 19080
rect 18340 19070 29400 19150
rect 6080 19060 29400 19070
rect 6080 18970 29400 18980
rect 6080 18960 18820 18970
rect 6080 18900 7270 18960
rect 7330 18900 18820 18960
rect 6080 18890 18820 18900
rect 18900 18890 29400 18970
rect 6080 18880 29400 18890
rect 6080 18700 29400 18800
<< metal4 >>
rect 3067 22490 3097 22576
rect 3343 22495 3373 22576
rect 3619 22495 3649 22576
rect 3895 22495 3925 22576
rect 4171 22495 4201 22576
rect 100 20245 300 22076
rect 100 20205 110 20245
rect 150 20205 170 20245
rect 210 20205 230 20245
rect 270 20205 300 20245
rect 100 500 300 20205
rect 400 21990 600 22076
rect 3060 22030 3105 22490
rect 3340 22035 3385 22495
rect 3615 22035 3660 22495
rect 3890 21990 3935 22495
rect 4170 21990 4210 22495
rect 4447 22490 4477 22576
rect 4445 22000 4485 22490
rect 4723 22485 4753 22576
rect 4999 22490 5029 22576
rect 4720 21995 4760 22485
rect 4995 22000 5035 22490
rect 5275 22485 5305 22576
rect 5551 22490 5581 22576
rect 5827 22490 5857 22576
rect 5270 21995 5310 22485
rect 5550 22000 5590 22490
rect 5825 22000 5865 22490
rect 6103 22485 6133 22576
rect 6379 22490 6409 22576
rect 6655 22490 6685 22576
rect 6931 22490 6961 22576
rect 7207 22490 7237 22576
rect 7483 22490 7513 22576
rect 7759 22490 7789 22576
rect 8035 22490 8065 22576
rect 8311 22490 8341 22576
rect 8587 22490 8617 22576
rect 8863 22490 8893 22576
rect 9139 22495 9169 22576
rect 9415 22495 9445 22576
rect 6100 21995 6140 22485
rect 6375 22000 6415 22490
rect 6650 22000 6690 22490
rect 6930 22000 6970 22490
rect 7205 22000 7245 22490
rect 7480 22040 7520 22490
rect 7755 22035 7795 22490
rect 8030 22035 8070 22490
rect 8310 22035 8350 22490
rect 8580 22030 8625 22490
rect 8860 22030 8905 22490
rect 9130 22030 9175 22495
rect 9410 22030 9455 22495
rect 9691 22476 9721 22576
rect 9967 22476 9997 22576
rect 10243 22476 10273 22576
rect 10519 22476 10549 22576
rect 10795 22476 10825 22576
rect 11071 22476 11101 22576
rect 11347 22476 11377 22576
rect 11623 22476 11653 22576
rect 11899 22490 11929 22576
rect 12175 22490 12205 22576
rect 12451 22570 12481 22576
rect 11895 22035 11940 22490
rect 400 21950 410 21990
rect 450 21950 470 21990
rect 510 21950 530 21990
rect 570 21950 600 21990
rect 400 19975 600 21950
rect 12175 21820 12215 22490
rect 12450 21900 12490 22570
rect 12727 22490 12757 22576
rect 13003 22490 13033 22576
rect 13279 22490 13309 22576
rect 13555 22490 13585 22576
rect 13831 22490 13861 22576
rect 12725 22030 12770 22490
rect 13000 22030 13045 22490
rect 13270 22030 13315 22490
rect 13550 22030 13595 22490
rect 13820 22030 13865 22490
rect 14107 22476 14137 22576
rect 14383 22476 14413 22576
rect 14659 22476 14689 22576
rect 400 19935 410 19975
rect 450 19935 470 19975
rect 510 19935 530 19975
rect 570 19935 600 19975
rect 400 500 600 19935
rect 6120 21840 6200 21928
rect 6680 21840 6750 21928
rect 7230 21840 7300 21928
rect 7780 21840 7850 21928
rect 8340 21840 8410 21928
rect 8890 21840 8960 21928
rect 9440 21840 9510 21928
rect 9990 21840 10060 21928
rect 10540 21840 10610 21928
rect 11100 21840 11170 21928
rect 11650 21840 11720 21928
rect 12200 21840 12270 21928
rect 12750 21840 12820 21934
rect 13300 21840 13370 21934
rect 13860 21840 13930 21934
rect 14410 21840 14480 21934
rect 6110 21830 6210 21840
rect 6110 21750 6130 21830
rect 6200 21750 6210 21830
rect 6110 21740 6210 21750
rect 6660 21830 6760 21840
rect 6660 21750 6680 21830
rect 6750 21750 6760 21830
rect 6660 21740 6760 21750
rect 7210 21830 7310 21840
rect 7210 21750 7230 21830
rect 7300 21750 7310 21830
rect 7210 21740 7310 21750
rect 7760 21830 7860 21840
rect 7760 21750 7780 21830
rect 7850 21750 7860 21830
rect 7760 21740 7860 21750
rect 8320 21830 8420 21840
rect 8320 21750 8340 21830
rect 8410 21750 8420 21830
rect 8320 21740 8420 21750
rect 8870 21830 8970 21840
rect 8870 21750 8890 21830
rect 8960 21750 8970 21830
rect 8870 21740 8970 21750
rect 9420 21830 9520 21840
rect 9420 21750 9440 21830
rect 9510 21750 9520 21830
rect 9420 21740 9520 21750
rect 9970 21830 10070 21840
rect 9970 21750 9990 21830
rect 10060 21750 10070 21830
rect 9970 21740 10070 21750
rect 10520 21830 10620 21840
rect 10520 21750 10540 21830
rect 10610 21750 10620 21830
rect 10520 21740 10620 21750
rect 11080 21830 11180 21840
rect 11080 21750 11100 21830
rect 11170 21750 11180 21830
rect 11080 21740 11180 21750
rect 11630 21830 11730 21840
rect 11630 21750 11650 21830
rect 11720 21750 11730 21830
rect 11630 21740 11730 21750
rect 12180 21830 12280 21840
rect 12180 21750 12200 21830
rect 12270 21750 12280 21830
rect 12180 21740 12280 21750
rect 12730 21830 12830 21840
rect 12730 21750 12750 21830
rect 12820 21750 12830 21830
rect 12730 21740 12830 21750
rect 13280 21830 13380 21840
rect 13280 21750 13300 21830
rect 13370 21750 13380 21830
rect 13280 21740 13380 21750
rect 13840 21830 13940 21840
rect 13840 21750 13860 21830
rect 13930 21750 13940 21830
rect 13840 21740 13940 21750
rect 14390 21830 14490 21840
rect 14390 21750 14410 21830
rect 14480 21750 14490 21830
rect 14390 21740 14490 21750
rect 14960 20240 15030 21934
rect 14950 20230 15040 20240
rect 14950 20150 14960 20230
rect 15030 20150 15040 20230
rect 14950 20140 15040 20150
rect 15510 20060 15580 21934
rect 15500 20050 15590 20060
rect 15500 19970 15510 20050
rect 15580 19970 15590 20050
rect 15500 19960 15590 19970
rect 16060 19880 16130 21934
rect 16050 19870 16140 19880
rect 16050 19790 16060 19870
rect 16130 19790 16140 19870
rect 16050 19780 16140 19790
rect 16620 19700 16690 21934
rect 16610 19690 16700 19700
rect 16610 19610 16620 19690
rect 16690 19610 16700 19690
rect 16610 19600 16700 19610
rect 17160 19520 17240 21934
rect 17150 19510 17250 19520
rect 17150 19430 17160 19510
rect 17240 19430 17250 19510
rect 17150 19420 17250 19430
rect 17720 19340 17800 21934
rect 17710 19330 17810 19340
rect 17710 19250 17720 19330
rect 17800 19250 17810 19330
rect 17710 19240 17810 19250
rect 18260 19160 18340 21934
rect 18250 19150 18350 19160
rect 18250 19070 18260 19150
rect 18340 19070 18350 19150
rect 18250 19060 18350 19070
rect 18820 18980 18900 21934
rect 23790 21660 23860 21934
rect 23770 21650 23870 21660
rect 23770 21570 23780 21650
rect 23860 21570 23870 21650
rect 23770 21560 23870 21570
rect 24350 21480 24410 21934
rect 24330 21470 24420 21480
rect 24330 21390 24340 21470
rect 24410 21390 24420 21470
rect 24330 21380 24420 21390
rect 24900 21310 24970 21934
rect 24870 21300 24990 21310
rect 24870 21220 24880 21300
rect 24980 21220 24990 21300
rect 24870 21210 24990 21220
rect 25450 21140 25530 21934
rect 25430 21130 25540 21140
rect 25430 21048 25450 21130
rect 25530 21048 25540 21130
rect 25430 21040 25540 21048
rect 26000 20960 26080 21934
rect 25980 20950 26090 20960
rect 25980 20870 26000 20950
rect 26080 20870 26090 20950
rect 25980 20860 26090 20870
rect 26540 20780 26620 21934
rect 26520 20770 26630 20780
rect 26520 20690 26540 20770
rect 26620 20690 26630 20770
rect 26520 20680 26630 20690
rect 27100 20600 27180 21934
rect 27080 20590 27190 20600
rect 27080 20510 27100 20590
rect 27180 20510 27190 20590
rect 27080 20500 27190 20510
rect 27640 20420 27720 21934
rect 27620 20410 27730 20420
rect 27620 20330 27640 20410
rect 27720 20330 27730 20410
rect 27620 20320 27730 20330
rect 18810 18970 18910 18980
rect 18810 18890 18820 18970
rect 18900 18890 18910 18970
rect 18810 18880 18910 18890
<< properties >>
string FIXED_BBOX 0 0 16100 22576
<< end >>
